magic
tech sky130A
magscale 1 2
timestamp 1623786739
<< obsli1 >>
rect 1104 1649 288880 287793
<< obsm1 >>
rect 290 688 289970 288108
<< metal2 >>
rect 1214 289200 1270 290000
rect 3698 289200 3754 290000
rect 6274 289200 6330 290000
rect 8758 289200 8814 290000
rect 11334 289200 11390 290000
rect 13910 289200 13966 290000
rect 16394 289200 16450 290000
rect 18970 289200 19026 290000
rect 21546 289200 21602 290000
rect 24030 289200 24086 290000
rect 26606 289200 26662 290000
rect 29182 289200 29238 290000
rect 31666 289200 31722 290000
rect 34242 289200 34298 290000
rect 36818 289200 36874 290000
rect 39302 289200 39358 290000
rect 41878 289200 41934 290000
rect 44454 289200 44510 290000
rect 46938 289200 46994 290000
rect 49514 289200 49570 290000
rect 51998 289200 52054 290000
rect 54574 289200 54630 290000
rect 57150 289200 57206 290000
rect 59634 289200 59690 290000
rect 62210 289200 62266 290000
rect 64786 289200 64842 290000
rect 67270 289200 67326 290000
rect 69846 289200 69902 290000
rect 72422 289200 72478 290000
rect 74906 289200 74962 290000
rect 77482 289200 77538 290000
rect 80058 289200 80114 290000
rect 82542 289200 82598 290000
rect 85118 289200 85174 290000
rect 87694 289200 87750 290000
rect 90178 289200 90234 290000
rect 92754 289200 92810 290000
rect 95330 289200 95386 290000
rect 97814 289200 97870 290000
rect 100390 289200 100446 290000
rect 102874 289200 102930 290000
rect 105450 289200 105506 290000
rect 108026 289200 108082 290000
rect 110510 289200 110566 290000
rect 113086 289200 113142 290000
rect 115662 289200 115718 290000
rect 118146 289200 118202 290000
rect 120722 289200 120778 290000
rect 123298 289200 123354 290000
rect 125782 289200 125838 290000
rect 128358 289200 128414 290000
rect 130934 289200 130990 290000
rect 133418 289200 133474 290000
rect 135994 289200 136050 290000
rect 138570 289200 138626 290000
rect 141054 289200 141110 290000
rect 143630 289200 143686 290000
rect 146206 289200 146262 290000
rect 148690 289200 148746 290000
rect 151266 289200 151322 290000
rect 153750 289200 153806 290000
rect 156326 289200 156382 290000
rect 158902 289200 158958 290000
rect 161386 289200 161442 290000
rect 163962 289200 164018 290000
rect 166538 289200 166594 290000
rect 169022 289200 169078 290000
rect 171598 289200 171654 290000
rect 174174 289200 174230 290000
rect 176658 289200 176714 290000
rect 179234 289200 179290 290000
rect 181810 289200 181866 290000
rect 184294 289200 184350 290000
rect 186870 289200 186926 290000
rect 189446 289200 189502 290000
rect 191930 289200 191986 290000
rect 194506 289200 194562 290000
rect 196990 289200 197046 290000
rect 199566 289200 199622 290000
rect 202142 289200 202198 290000
rect 204626 289200 204682 290000
rect 207202 289200 207258 290000
rect 209778 289200 209834 290000
rect 212262 289200 212318 290000
rect 214838 289200 214894 290000
rect 217414 289200 217470 290000
rect 219898 289200 219954 290000
rect 222474 289200 222530 290000
rect 225050 289200 225106 290000
rect 227534 289200 227590 290000
rect 230110 289200 230166 290000
rect 232686 289200 232742 290000
rect 235170 289200 235226 290000
rect 237746 289200 237802 290000
rect 240322 289200 240378 290000
rect 242806 289200 242862 290000
rect 245382 289200 245438 290000
rect 247866 289200 247922 290000
rect 250442 289200 250498 290000
rect 253018 289200 253074 290000
rect 255502 289200 255558 290000
rect 258078 289200 258134 290000
rect 260654 289200 260710 290000
rect 263138 289200 263194 290000
rect 265714 289200 265770 290000
rect 268290 289200 268346 290000
rect 270774 289200 270830 290000
rect 273350 289200 273406 290000
rect 275926 289200 275982 290000
rect 278410 289200 278466 290000
rect 280986 289200 281042 290000
rect 283562 289200 283618 290000
rect 286046 289200 286102 290000
rect 288622 289200 288678 290000
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 2042 0 2098 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3790 0 3846 800
rect 4342 0 4398 800
rect 4986 0 5042 800
rect 5538 0 5594 800
rect 6182 0 6238 800
rect 6734 0 6790 800
rect 7378 0 7434 800
rect 7930 0 7986 800
rect 8482 0 8538 800
rect 9126 0 9182 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11426 0 11482 800
rect 12070 0 12126 800
rect 12622 0 12678 800
rect 13266 0 13322 800
rect 13818 0 13874 800
rect 14462 0 14518 800
rect 15014 0 15070 800
rect 15566 0 15622 800
rect 16210 0 16266 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 17958 0 18014 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20350 0 20406 800
rect 20902 0 20958 800
rect 21546 0 21602 800
rect 22098 0 22154 800
rect 22650 0 22706 800
rect 23294 0 23350 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25042 0 25098 800
rect 25686 0 25742 800
rect 26238 0 26294 800
rect 26790 0 26846 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28630 0 28686 800
rect 29182 0 29238 800
rect 29734 0 29790 800
rect 30378 0 30434 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32126 0 32182 800
rect 32770 0 32826 800
rect 33322 0 33378 800
rect 33874 0 33930 800
rect 34518 0 34574 800
rect 35070 0 35126 800
rect 35714 0 35770 800
rect 36266 0 36322 800
rect 36910 0 36966 800
rect 37462 0 37518 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39210 0 39266 800
rect 39854 0 39910 800
rect 40406 0 40462 800
rect 40958 0 41014 800
rect 41602 0 41658 800
rect 42154 0 42210 800
rect 42798 0 42854 800
rect 43350 0 43406 800
rect 43994 0 44050 800
rect 44546 0 44602 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 46294 0 46350 800
rect 46938 0 46994 800
rect 47490 0 47546 800
rect 48042 0 48098 800
rect 48686 0 48742 800
rect 49238 0 49294 800
rect 49882 0 49938 800
rect 50434 0 50490 800
rect 51078 0 51134 800
rect 51630 0 51686 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 53378 0 53434 800
rect 54022 0 54078 800
rect 54574 0 54630 800
rect 55218 0 55274 800
rect 55770 0 55826 800
rect 56322 0 56378 800
rect 56966 0 57022 800
rect 57518 0 57574 800
rect 58162 0 58218 800
rect 58714 0 58770 800
rect 59266 0 59322 800
rect 59910 0 59966 800
rect 60462 0 60518 800
rect 61106 0 61162 800
rect 61658 0 61714 800
rect 62302 0 62358 800
rect 62854 0 62910 800
rect 63406 0 63462 800
rect 64050 0 64106 800
rect 64602 0 64658 800
rect 65246 0 65302 800
rect 65798 0 65854 800
rect 66350 0 66406 800
rect 66994 0 67050 800
rect 67546 0 67602 800
rect 68190 0 68246 800
rect 68742 0 68798 800
rect 69386 0 69442 800
rect 69938 0 69994 800
rect 70490 0 70546 800
rect 71134 0 71190 800
rect 71686 0 71742 800
rect 72330 0 72386 800
rect 72882 0 72938 800
rect 73526 0 73582 800
rect 74078 0 74134 800
rect 74630 0 74686 800
rect 75274 0 75330 800
rect 75826 0 75882 800
rect 76470 0 76526 800
rect 77022 0 77078 800
rect 77574 0 77630 800
rect 78218 0 78274 800
rect 78770 0 78826 800
rect 79414 0 79470 800
rect 79966 0 80022 800
rect 80610 0 80666 800
rect 81162 0 81218 800
rect 81714 0 81770 800
rect 82358 0 82414 800
rect 82910 0 82966 800
rect 83554 0 83610 800
rect 84106 0 84162 800
rect 84658 0 84714 800
rect 85302 0 85358 800
rect 85854 0 85910 800
rect 86498 0 86554 800
rect 87050 0 87106 800
rect 87694 0 87750 800
rect 88246 0 88302 800
rect 88798 0 88854 800
rect 89442 0 89498 800
rect 89994 0 90050 800
rect 90638 0 90694 800
rect 91190 0 91246 800
rect 91834 0 91890 800
rect 92386 0 92442 800
rect 92938 0 92994 800
rect 93582 0 93638 800
rect 94134 0 94190 800
rect 94778 0 94834 800
rect 95330 0 95386 800
rect 95882 0 95938 800
rect 96526 0 96582 800
rect 97078 0 97134 800
rect 97722 0 97778 800
rect 98274 0 98330 800
rect 98918 0 98974 800
rect 99470 0 99526 800
rect 100022 0 100078 800
rect 100666 0 100722 800
rect 101218 0 101274 800
rect 101862 0 101918 800
rect 102414 0 102470 800
rect 103058 0 103114 800
rect 103610 0 103666 800
rect 104162 0 104218 800
rect 104806 0 104862 800
rect 105358 0 105414 800
rect 106002 0 106058 800
rect 106554 0 106610 800
rect 107106 0 107162 800
rect 107750 0 107806 800
rect 108302 0 108358 800
rect 108946 0 109002 800
rect 109498 0 109554 800
rect 110142 0 110198 800
rect 110694 0 110750 800
rect 111246 0 111302 800
rect 111890 0 111946 800
rect 112442 0 112498 800
rect 113086 0 113142 800
rect 113638 0 113694 800
rect 114190 0 114246 800
rect 114834 0 114890 800
rect 115386 0 115442 800
rect 116030 0 116086 800
rect 116582 0 116638 800
rect 117226 0 117282 800
rect 117778 0 117834 800
rect 118330 0 118386 800
rect 118974 0 119030 800
rect 119526 0 119582 800
rect 120170 0 120226 800
rect 120722 0 120778 800
rect 121366 0 121422 800
rect 121918 0 121974 800
rect 122470 0 122526 800
rect 123114 0 123170 800
rect 123666 0 123722 800
rect 124310 0 124366 800
rect 124862 0 124918 800
rect 125414 0 125470 800
rect 126058 0 126114 800
rect 126610 0 126666 800
rect 127254 0 127310 800
rect 127806 0 127862 800
rect 128450 0 128506 800
rect 129002 0 129058 800
rect 129554 0 129610 800
rect 130198 0 130254 800
rect 130750 0 130806 800
rect 131394 0 131450 800
rect 131946 0 132002 800
rect 132498 0 132554 800
rect 133142 0 133198 800
rect 133694 0 133750 800
rect 134338 0 134394 800
rect 134890 0 134946 800
rect 135534 0 135590 800
rect 136086 0 136142 800
rect 136638 0 136694 800
rect 137282 0 137338 800
rect 137834 0 137890 800
rect 138478 0 138534 800
rect 139030 0 139086 800
rect 139674 0 139730 800
rect 140226 0 140282 800
rect 140778 0 140834 800
rect 141422 0 141478 800
rect 141974 0 142030 800
rect 142618 0 142674 800
rect 143170 0 143226 800
rect 143722 0 143778 800
rect 144366 0 144422 800
rect 144918 0 144974 800
rect 145562 0 145618 800
rect 146114 0 146170 800
rect 146758 0 146814 800
rect 147310 0 147366 800
rect 147862 0 147918 800
rect 148506 0 148562 800
rect 149058 0 149114 800
rect 149702 0 149758 800
rect 150254 0 150310 800
rect 150806 0 150862 800
rect 151450 0 151506 800
rect 152002 0 152058 800
rect 152646 0 152702 800
rect 153198 0 153254 800
rect 153842 0 153898 800
rect 154394 0 154450 800
rect 154946 0 155002 800
rect 155590 0 155646 800
rect 156142 0 156198 800
rect 156786 0 156842 800
rect 157338 0 157394 800
rect 157982 0 158038 800
rect 158534 0 158590 800
rect 159086 0 159142 800
rect 159730 0 159786 800
rect 160282 0 160338 800
rect 160926 0 160982 800
rect 161478 0 161534 800
rect 162030 0 162086 800
rect 162674 0 162730 800
rect 163226 0 163282 800
rect 163870 0 163926 800
rect 164422 0 164478 800
rect 165066 0 165122 800
rect 165618 0 165674 800
rect 166170 0 166226 800
rect 166814 0 166870 800
rect 167366 0 167422 800
rect 168010 0 168066 800
rect 168562 0 168618 800
rect 169114 0 169170 800
rect 169758 0 169814 800
rect 170310 0 170366 800
rect 170954 0 171010 800
rect 171506 0 171562 800
rect 172150 0 172206 800
rect 172702 0 172758 800
rect 173254 0 173310 800
rect 173898 0 173954 800
rect 174450 0 174506 800
rect 175094 0 175150 800
rect 175646 0 175702 800
rect 176290 0 176346 800
rect 176842 0 176898 800
rect 177394 0 177450 800
rect 178038 0 178094 800
rect 178590 0 178646 800
rect 179234 0 179290 800
rect 179786 0 179842 800
rect 180338 0 180394 800
rect 180982 0 181038 800
rect 181534 0 181590 800
rect 182178 0 182234 800
rect 182730 0 182786 800
rect 183374 0 183430 800
rect 183926 0 183982 800
rect 184478 0 184534 800
rect 185122 0 185178 800
rect 185674 0 185730 800
rect 186318 0 186374 800
rect 186870 0 186926 800
rect 187422 0 187478 800
rect 188066 0 188122 800
rect 188618 0 188674 800
rect 189262 0 189318 800
rect 189814 0 189870 800
rect 190458 0 190514 800
rect 191010 0 191066 800
rect 191562 0 191618 800
rect 192206 0 192262 800
rect 192758 0 192814 800
rect 193402 0 193458 800
rect 193954 0 194010 800
rect 194598 0 194654 800
rect 195150 0 195206 800
rect 195702 0 195758 800
rect 196346 0 196402 800
rect 196898 0 196954 800
rect 197542 0 197598 800
rect 198094 0 198150 800
rect 198646 0 198702 800
rect 199290 0 199346 800
rect 199842 0 199898 800
rect 200486 0 200542 800
rect 201038 0 201094 800
rect 201682 0 201738 800
rect 202234 0 202290 800
rect 202786 0 202842 800
rect 203430 0 203486 800
rect 203982 0 204038 800
rect 204626 0 204682 800
rect 205178 0 205234 800
rect 205822 0 205878 800
rect 206374 0 206430 800
rect 206926 0 206982 800
rect 207570 0 207626 800
rect 208122 0 208178 800
rect 208766 0 208822 800
rect 209318 0 209374 800
rect 209870 0 209926 800
rect 210514 0 210570 800
rect 211066 0 211122 800
rect 211710 0 211766 800
rect 212262 0 212318 800
rect 212906 0 212962 800
rect 213458 0 213514 800
rect 214010 0 214066 800
rect 214654 0 214710 800
rect 215206 0 215262 800
rect 215850 0 215906 800
rect 216402 0 216458 800
rect 216954 0 217010 800
rect 217598 0 217654 800
rect 218150 0 218206 800
rect 218794 0 218850 800
rect 219346 0 219402 800
rect 219990 0 220046 800
rect 220542 0 220598 800
rect 221094 0 221150 800
rect 221738 0 221794 800
rect 222290 0 222346 800
rect 222934 0 222990 800
rect 223486 0 223542 800
rect 224130 0 224186 800
rect 224682 0 224738 800
rect 225234 0 225290 800
rect 225878 0 225934 800
rect 226430 0 226486 800
rect 227074 0 227130 800
rect 227626 0 227682 800
rect 228178 0 228234 800
rect 228822 0 228878 800
rect 229374 0 229430 800
rect 230018 0 230074 800
rect 230570 0 230626 800
rect 231214 0 231270 800
rect 231766 0 231822 800
rect 232318 0 232374 800
rect 232962 0 233018 800
rect 233514 0 233570 800
rect 234158 0 234214 800
rect 234710 0 234766 800
rect 235262 0 235318 800
rect 235906 0 235962 800
rect 236458 0 236514 800
rect 237102 0 237158 800
rect 237654 0 237710 800
rect 238298 0 238354 800
rect 238850 0 238906 800
rect 239402 0 239458 800
rect 240046 0 240102 800
rect 240598 0 240654 800
rect 241242 0 241298 800
rect 241794 0 241850 800
rect 242438 0 242494 800
rect 242990 0 243046 800
rect 243542 0 243598 800
rect 244186 0 244242 800
rect 244738 0 244794 800
rect 245382 0 245438 800
rect 245934 0 245990 800
rect 246486 0 246542 800
rect 247130 0 247186 800
rect 247682 0 247738 800
rect 248326 0 248382 800
rect 248878 0 248934 800
rect 249522 0 249578 800
rect 250074 0 250130 800
rect 250626 0 250682 800
rect 251270 0 251326 800
rect 251822 0 251878 800
rect 252466 0 252522 800
rect 253018 0 253074 800
rect 253570 0 253626 800
rect 254214 0 254270 800
rect 254766 0 254822 800
rect 255410 0 255466 800
rect 255962 0 256018 800
rect 256606 0 256662 800
rect 257158 0 257214 800
rect 257710 0 257766 800
rect 258354 0 258410 800
rect 258906 0 258962 800
rect 259550 0 259606 800
rect 260102 0 260158 800
rect 260746 0 260802 800
rect 261298 0 261354 800
rect 261850 0 261906 800
rect 262494 0 262550 800
rect 263046 0 263102 800
rect 263690 0 263746 800
rect 264242 0 264298 800
rect 264794 0 264850 800
rect 265438 0 265494 800
rect 265990 0 266046 800
rect 266634 0 266690 800
rect 267186 0 267242 800
rect 267830 0 267886 800
rect 268382 0 268438 800
rect 268934 0 268990 800
rect 269578 0 269634 800
rect 270130 0 270186 800
rect 270774 0 270830 800
rect 271326 0 271382 800
rect 271878 0 271934 800
rect 272522 0 272578 800
rect 273074 0 273130 800
rect 273718 0 273774 800
rect 274270 0 274326 800
rect 274914 0 274970 800
rect 275466 0 275522 800
rect 276018 0 276074 800
rect 276662 0 276718 800
rect 277214 0 277270 800
rect 277858 0 277914 800
rect 278410 0 278466 800
rect 279054 0 279110 800
rect 279606 0 279662 800
rect 280158 0 280214 800
rect 280802 0 280858 800
rect 281354 0 281410 800
rect 281998 0 282054 800
rect 282550 0 282606 800
rect 283102 0 283158 800
rect 283746 0 283802 800
rect 284298 0 284354 800
rect 284942 0 284998 800
rect 285494 0 285550 800
rect 286138 0 286194 800
rect 286690 0 286746 800
rect 287242 0 287298 800
rect 287886 0 287942 800
rect 288438 0 288494 800
rect 289082 0 289138 800
rect 289634 0 289690 800
<< obsm2 >>
rect 296 289144 1158 289200
rect 1326 289144 3642 289200
rect 3810 289144 6218 289200
rect 6386 289144 8702 289200
rect 8870 289144 11278 289200
rect 11446 289144 13854 289200
rect 14022 289144 16338 289200
rect 16506 289144 18914 289200
rect 19082 289144 21490 289200
rect 21658 289144 23974 289200
rect 24142 289144 26550 289200
rect 26718 289144 29126 289200
rect 29294 289144 31610 289200
rect 31778 289144 34186 289200
rect 34354 289144 36762 289200
rect 36930 289144 39246 289200
rect 39414 289144 41822 289200
rect 41990 289144 44398 289200
rect 44566 289144 46882 289200
rect 47050 289144 49458 289200
rect 49626 289144 51942 289200
rect 52110 289144 54518 289200
rect 54686 289144 57094 289200
rect 57262 289144 59578 289200
rect 59746 289144 62154 289200
rect 62322 289144 64730 289200
rect 64898 289144 67214 289200
rect 67382 289144 69790 289200
rect 69958 289144 72366 289200
rect 72534 289144 74850 289200
rect 75018 289144 77426 289200
rect 77594 289144 80002 289200
rect 80170 289144 82486 289200
rect 82654 289144 85062 289200
rect 85230 289144 87638 289200
rect 87806 289144 90122 289200
rect 90290 289144 92698 289200
rect 92866 289144 95274 289200
rect 95442 289144 97758 289200
rect 97926 289144 100334 289200
rect 100502 289144 102818 289200
rect 102986 289144 105394 289200
rect 105562 289144 107970 289200
rect 108138 289144 110454 289200
rect 110622 289144 113030 289200
rect 113198 289144 115606 289200
rect 115774 289144 118090 289200
rect 118258 289144 120666 289200
rect 120834 289144 123242 289200
rect 123410 289144 125726 289200
rect 125894 289144 128302 289200
rect 128470 289144 130878 289200
rect 131046 289144 133362 289200
rect 133530 289144 135938 289200
rect 136106 289144 138514 289200
rect 138682 289144 140998 289200
rect 141166 289144 143574 289200
rect 143742 289144 146150 289200
rect 146318 289144 148634 289200
rect 148802 289144 151210 289200
rect 151378 289144 153694 289200
rect 153862 289144 156270 289200
rect 156438 289144 158846 289200
rect 159014 289144 161330 289200
rect 161498 289144 163906 289200
rect 164074 289144 166482 289200
rect 166650 289144 168966 289200
rect 169134 289144 171542 289200
rect 171710 289144 174118 289200
rect 174286 289144 176602 289200
rect 176770 289144 179178 289200
rect 179346 289144 181754 289200
rect 181922 289144 184238 289200
rect 184406 289144 186814 289200
rect 186982 289144 189390 289200
rect 189558 289144 191874 289200
rect 192042 289144 194450 289200
rect 194618 289144 196934 289200
rect 197102 289144 199510 289200
rect 199678 289144 202086 289200
rect 202254 289144 204570 289200
rect 204738 289144 207146 289200
rect 207314 289144 209722 289200
rect 209890 289144 212206 289200
rect 212374 289144 214782 289200
rect 214950 289144 217358 289200
rect 217526 289144 219842 289200
rect 220010 289144 222418 289200
rect 222586 289144 224994 289200
rect 225162 289144 227478 289200
rect 227646 289144 230054 289200
rect 230222 289144 232630 289200
rect 232798 289144 235114 289200
rect 235282 289144 237690 289200
rect 237858 289144 240266 289200
rect 240434 289144 242750 289200
rect 242918 289144 245326 289200
rect 245494 289144 247810 289200
rect 247978 289144 250386 289200
rect 250554 289144 252962 289200
rect 253130 289144 255446 289200
rect 255614 289144 258022 289200
rect 258190 289144 260598 289200
rect 260766 289144 263082 289200
rect 263250 289144 265658 289200
rect 265826 289144 268234 289200
rect 268402 289144 270718 289200
rect 270886 289144 273294 289200
rect 273462 289144 275870 289200
rect 276038 289144 278354 289200
rect 278522 289144 280930 289200
rect 281098 289144 283506 289200
rect 283674 289144 285990 289200
rect 286158 289144 288566 289200
rect 288734 289144 289966 289200
rect 296 856 289966 289144
rect 406 682 790 856
rect 958 682 1342 856
rect 1510 682 1986 856
rect 2154 682 2538 856
rect 2706 682 3182 856
rect 3350 682 3734 856
rect 3902 682 4286 856
rect 4454 682 4930 856
rect 5098 682 5482 856
rect 5650 682 6126 856
rect 6294 682 6678 856
rect 6846 682 7322 856
rect 7490 682 7874 856
rect 8042 682 8426 856
rect 8594 682 9070 856
rect 9238 682 9622 856
rect 9790 682 10266 856
rect 10434 682 10818 856
rect 10986 682 11370 856
rect 11538 682 12014 856
rect 12182 682 12566 856
rect 12734 682 13210 856
rect 13378 682 13762 856
rect 13930 682 14406 856
rect 14574 682 14958 856
rect 15126 682 15510 856
rect 15678 682 16154 856
rect 16322 682 16706 856
rect 16874 682 17350 856
rect 17518 682 17902 856
rect 18070 682 18546 856
rect 18714 682 19098 856
rect 19266 682 19650 856
rect 19818 682 20294 856
rect 20462 682 20846 856
rect 21014 682 21490 856
rect 21658 682 22042 856
rect 22210 682 22594 856
rect 22762 682 23238 856
rect 23406 682 23790 856
rect 23958 682 24434 856
rect 24602 682 24986 856
rect 25154 682 25630 856
rect 25798 682 26182 856
rect 26350 682 26734 856
rect 26902 682 27378 856
rect 27546 682 27930 856
rect 28098 682 28574 856
rect 28742 682 29126 856
rect 29294 682 29678 856
rect 29846 682 30322 856
rect 30490 682 30874 856
rect 31042 682 31518 856
rect 31686 682 32070 856
rect 32238 682 32714 856
rect 32882 682 33266 856
rect 33434 682 33818 856
rect 33986 682 34462 856
rect 34630 682 35014 856
rect 35182 682 35658 856
rect 35826 682 36210 856
rect 36378 682 36854 856
rect 37022 682 37406 856
rect 37574 682 37958 856
rect 38126 682 38602 856
rect 38770 682 39154 856
rect 39322 682 39798 856
rect 39966 682 40350 856
rect 40518 682 40902 856
rect 41070 682 41546 856
rect 41714 682 42098 856
rect 42266 682 42742 856
rect 42910 682 43294 856
rect 43462 682 43938 856
rect 44106 682 44490 856
rect 44658 682 45042 856
rect 45210 682 45686 856
rect 45854 682 46238 856
rect 46406 682 46882 856
rect 47050 682 47434 856
rect 47602 682 47986 856
rect 48154 682 48630 856
rect 48798 682 49182 856
rect 49350 682 49826 856
rect 49994 682 50378 856
rect 50546 682 51022 856
rect 51190 682 51574 856
rect 51742 682 52126 856
rect 52294 682 52770 856
rect 52938 682 53322 856
rect 53490 682 53966 856
rect 54134 682 54518 856
rect 54686 682 55162 856
rect 55330 682 55714 856
rect 55882 682 56266 856
rect 56434 682 56910 856
rect 57078 682 57462 856
rect 57630 682 58106 856
rect 58274 682 58658 856
rect 58826 682 59210 856
rect 59378 682 59854 856
rect 60022 682 60406 856
rect 60574 682 61050 856
rect 61218 682 61602 856
rect 61770 682 62246 856
rect 62414 682 62798 856
rect 62966 682 63350 856
rect 63518 682 63994 856
rect 64162 682 64546 856
rect 64714 682 65190 856
rect 65358 682 65742 856
rect 65910 682 66294 856
rect 66462 682 66938 856
rect 67106 682 67490 856
rect 67658 682 68134 856
rect 68302 682 68686 856
rect 68854 682 69330 856
rect 69498 682 69882 856
rect 70050 682 70434 856
rect 70602 682 71078 856
rect 71246 682 71630 856
rect 71798 682 72274 856
rect 72442 682 72826 856
rect 72994 682 73470 856
rect 73638 682 74022 856
rect 74190 682 74574 856
rect 74742 682 75218 856
rect 75386 682 75770 856
rect 75938 682 76414 856
rect 76582 682 76966 856
rect 77134 682 77518 856
rect 77686 682 78162 856
rect 78330 682 78714 856
rect 78882 682 79358 856
rect 79526 682 79910 856
rect 80078 682 80554 856
rect 80722 682 81106 856
rect 81274 682 81658 856
rect 81826 682 82302 856
rect 82470 682 82854 856
rect 83022 682 83498 856
rect 83666 682 84050 856
rect 84218 682 84602 856
rect 84770 682 85246 856
rect 85414 682 85798 856
rect 85966 682 86442 856
rect 86610 682 86994 856
rect 87162 682 87638 856
rect 87806 682 88190 856
rect 88358 682 88742 856
rect 88910 682 89386 856
rect 89554 682 89938 856
rect 90106 682 90582 856
rect 90750 682 91134 856
rect 91302 682 91778 856
rect 91946 682 92330 856
rect 92498 682 92882 856
rect 93050 682 93526 856
rect 93694 682 94078 856
rect 94246 682 94722 856
rect 94890 682 95274 856
rect 95442 682 95826 856
rect 95994 682 96470 856
rect 96638 682 97022 856
rect 97190 682 97666 856
rect 97834 682 98218 856
rect 98386 682 98862 856
rect 99030 682 99414 856
rect 99582 682 99966 856
rect 100134 682 100610 856
rect 100778 682 101162 856
rect 101330 682 101806 856
rect 101974 682 102358 856
rect 102526 682 103002 856
rect 103170 682 103554 856
rect 103722 682 104106 856
rect 104274 682 104750 856
rect 104918 682 105302 856
rect 105470 682 105946 856
rect 106114 682 106498 856
rect 106666 682 107050 856
rect 107218 682 107694 856
rect 107862 682 108246 856
rect 108414 682 108890 856
rect 109058 682 109442 856
rect 109610 682 110086 856
rect 110254 682 110638 856
rect 110806 682 111190 856
rect 111358 682 111834 856
rect 112002 682 112386 856
rect 112554 682 113030 856
rect 113198 682 113582 856
rect 113750 682 114134 856
rect 114302 682 114778 856
rect 114946 682 115330 856
rect 115498 682 115974 856
rect 116142 682 116526 856
rect 116694 682 117170 856
rect 117338 682 117722 856
rect 117890 682 118274 856
rect 118442 682 118918 856
rect 119086 682 119470 856
rect 119638 682 120114 856
rect 120282 682 120666 856
rect 120834 682 121310 856
rect 121478 682 121862 856
rect 122030 682 122414 856
rect 122582 682 123058 856
rect 123226 682 123610 856
rect 123778 682 124254 856
rect 124422 682 124806 856
rect 124974 682 125358 856
rect 125526 682 126002 856
rect 126170 682 126554 856
rect 126722 682 127198 856
rect 127366 682 127750 856
rect 127918 682 128394 856
rect 128562 682 128946 856
rect 129114 682 129498 856
rect 129666 682 130142 856
rect 130310 682 130694 856
rect 130862 682 131338 856
rect 131506 682 131890 856
rect 132058 682 132442 856
rect 132610 682 133086 856
rect 133254 682 133638 856
rect 133806 682 134282 856
rect 134450 682 134834 856
rect 135002 682 135478 856
rect 135646 682 136030 856
rect 136198 682 136582 856
rect 136750 682 137226 856
rect 137394 682 137778 856
rect 137946 682 138422 856
rect 138590 682 138974 856
rect 139142 682 139618 856
rect 139786 682 140170 856
rect 140338 682 140722 856
rect 140890 682 141366 856
rect 141534 682 141918 856
rect 142086 682 142562 856
rect 142730 682 143114 856
rect 143282 682 143666 856
rect 143834 682 144310 856
rect 144478 682 144862 856
rect 145030 682 145506 856
rect 145674 682 146058 856
rect 146226 682 146702 856
rect 146870 682 147254 856
rect 147422 682 147806 856
rect 147974 682 148450 856
rect 148618 682 149002 856
rect 149170 682 149646 856
rect 149814 682 150198 856
rect 150366 682 150750 856
rect 150918 682 151394 856
rect 151562 682 151946 856
rect 152114 682 152590 856
rect 152758 682 153142 856
rect 153310 682 153786 856
rect 153954 682 154338 856
rect 154506 682 154890 856
rect 155058 682 155534 856
rect 155702 682 156086 856
rect 156254 682 156730 856
rect 156898 682 157282 856
rect 157450 682 157926 856
rect 158094 682 158478 856
rect 158646 682 159030 856
rect 159198 682 159674 856
rect 159842 682 160226 856
rect 160394 682 160870 856
rect 161038 682 161422 856
rect 161590 682 161974 856
rect 162142 682 162618 856
rect 162786 682 163170 856
rect 163338 682 163814 856
rect 163982 682 164366 856
rect 164534 682 165010 856
rect 165178 682 165562 856
rect 165730 682 166114 856
rect 166282 682 166758 856
rect 166926 682 167310 856
rect 167478 682 167954 856
rect 168122 682 168506 856
rect 168674 682 169058 856
rect 169226 682 169702 856
rect 169870 682 170254 856
rect 170422 682 170898 856
rect 171066 682 171450 856
rect 171618 682 172094 856
rect 172262 682 172646 856
rect 172814 682 173198 856
rect 173366 682 173842 856
rect 174010 682 174394 856
rect 174562 682 175038 856
rect 175206 682 175590 856
rect 175758 682 176234 856
rect 176402 682 176786 856
rect 176954 682 177338 856
rect 177506 682 177982 856
rect 178150 682 178534 856
rect 178702 682 179178 856
rect 179346 682 179730 856
rect 179898 682 180282 856
rect 180450 682 180926 856
rect 181094 682 181478 856
rect 181646 682 182122 856
rect 182290 682 182674 856
rect 182842 682 183318 856
rect 183486 682 183870 856
rect 184038 682 184422 856
rect 184590 682 185066 856
rect 185234 682 185618 856
rect 185786 682 186262 856
rect 186430 682 186814 856
rect 186982 682 187366 856
rect 187534 682 188010 856
rect 188178 682 188562 856
rect 188730 682 189206 856
rect 189374 682 189758 856
rect 189926 682 190402 856
rect 190570 682 190954 856
rect 191122 682 191506 856
rect 191674 682 192150 856
rect 192318 682 192702 856
rect 192870 682 193346 856
rect 193514 682 193898 856
rect 194066 682 194542 856
rect 194710 682 195094 856
rect 195262 682 195646 856
rect 195814 682 196290 856
rect 196458 682 196842 856
rect 197010 682 197486 856
rect 197654 682 198038 856
rect 198206 682 198590 856
rect 198758 682 199234 856
rect 199402 682 199786 856
rect 199954 682 200430 856
rect 200598 682 200982 856
rect 201150 682 201626 856
rect 201794 682 202178 856
rect 202346 682 202730 856
rect 202898 682 203374 856
rect 203542 682 203926 856
rect 204094 682 204570 856
rect 204738 682 205122 856
rect 205290 682 205766 856
rect 205934 682 206318 856
rect 206486 682 206870 856
rect 207038 682 207514 856
rect 207682 682 208066 856
rect 208234 682 208710 856
rect 208878 682 209262 856
rect 209430 682 209814 856
rect 209982 682 210458 856
rect 210626 682 211010 856
rect 211178 682 211654 856
rect 211822 682 212206 856
rect 212374 682 212850 856
rect 213018 682 213402 856
rect 213570 682 213954 856
rect 214122 682 214598 856
rect 214766 682 215150 856
rect 215318 682 215794 856
rect 215962 682 216346 856
rect 216514 682 216898 856
rect 217066 682 217542 856
rect 217710 682 218094 856
rect 218262 682 218738 856
rect 218906 682 219290 856
rect 219458 682 219934 856
rect 220102 682 220486 856
rect 220654 682 221038 856
rect 221206 682 221682 856
rect 221850 682 222234 856
rect 222402 682 222878 856
rect 223046 682 223430 856
rect 223598 682 224074 856
rect 224242 682 224626 856
rect 224794 682 225178 856
rect 225346 682 225822 856
rect 225990 682 226374 856
rect 226542 682 227018 856
rect 227186 682 227570 856
rect 227738 682 228122 856
rect 228290 682 228766 856
rect 228934 682 229318 856
rect 229486 682 229962 856
rect 230130 682 230514 856
rect 230682 682 231158 856
rect 231326 682 231710 856
rect 231878 682 232262 856
rect 232430 682 232906 856
rect 233074 682 233458 856
rect 233626 682 234102 856
rect 234270 682 234654 856
rect 234822 682 235206 856
rect 235374 682 235850 856
rect 236018 682 236402 856
rect 236570 682 237046 856
rect 237214 682 237598 856
rect 237766 682 238242 856
rect 238410 682 238794 856
rect 238962 682 239346 856
rect 239514 682 239990 856
rect 240158 682 240542 856
rect 240710 682 241186 856
rect 241354 682 241738 856
rect 241906 682 242382 856
rect 242550 682 242934 856
rect 243102 682 243486 856
rect 243654 682 244130 856
rect 244298 682 244682 856
rect 244850 682 245326 856
rect 245494 682 245878 856
rect 246046 682 246430 856
rect 246598 682 247074 856
rect 247242 682 247626 856
rect 247794 682 248270 856
rect 248438 682 248822 856
rect 248990 682 249466 856
rect 249634 682 250018 856
rect 250186 682 250570 856
rect 250738 682 251214 856
rect 251382 682 251766 856
rect 251934 682 252410 856
rect 252578 682 252962 856
rect 253130 682 253514 856
rect 253682 682 254158 856
rect 254326 682 254710 856
rect 254878 682 255354 856
rect 255522 682 255906 856
rect 256074 682 256550 856
rect 256718 682 257102 856
rect 257270 682 257654 856
rect 257822 682 258298 856
rect 258466 682 258850 856
rect 259018 682 259494 856
rect 259662 682 260046 856
rect 260214 682 260690 856
rect 260858 682 261242 856
rect 261410 682 261794 856
rect 261962 682 262438 856
rect 262606 682 262990 856
rect 263158 682 263634 856
rect 263802 682 264186 856
rect 264354 682 264738 856
rect 264906 682 265382 856
rect 265550 682 265934 856
rect 266102 682 266578 856
rect 266746 682 267130 856
rect 267298 682 267774 856
rect 267942 682 268326 856
rect 268494 682 268878 856
rect 269046 682 269522 856
rect 269690 682 270074 856
rect 270242 682 270718 856
rect 270886 682 271270 856
rect 271438 682 271822 856
rect 271990 682 272466 856
rect 272634 682 273018 856
rect 273186 682 273662 856
rect 273830 682 274214 856
rect 274382 682 274858 856
rect 275026 682 275410 856
rect 275578 682 275962 856
rect 276130 682 276606 856
rect 276774 682 277158 856
rect 277326 682 277802 856
rect 277970 682 278354 856
rect 278522 682 278998 856
rect 279166 682 279550 856
rect 279718 682 280102 856
rect 280270 682 280746 856
rect 280914 682 281298 856
rect 281466 682 281942 856
rect 282110 682 282494 856
rect 282662 682 283046 856
rect 283214 682 283690 856
rect 283858 682 284242 856
rect 284410 682 284886 856
rect 285054 682 285438 856
rect 285606 682 286082 856
rect 286250 682 286634 856
rect 286802 682 287186 856
rect 287354 682 287830 856
rect 287998 682 288382 856
rect 288550 682 289026 856
rect 289194 682 289578 856
rect 289746 682 289966 856
<< metal3 >>
rect 289200 217472 290000 217592
rect 0 144984 800 145104
rect 289200 72496 290000 72616
<< obsm3 >>
rect 800 217672 289971 287809
rect 800 217392 289120 217672
rect 800 145184 289971 217392
rect 880 144904 289971 145184
rect 800 72696 289971 144904
rect 800 72416 289120 72696
rect 800 1259 289971 72416
<< metal4 >>
rect 4208 2128 4528 287824
rect 4868 2176 5188 287776
rect 5528 2176 5848 287776
rect 6188 2176 6508 287776
rect 19568 2128 19888 287824
rect 20228 2176 20548 287776
rect 20888 2176 21208 287776
rect 21548 2176 21868 287776
rect 34928 2128 35248 287824
rect 35588 2176 35908 287776
rect 36248 2176 36568 287776
rect 36908 2176 37228 287776
rect 50288 2128 50608 287824
rect 50948 2176 51268 287776
rect 51608 2176 51928 287776
rect 52268 2176 52588 287776
rect 65648 2128 65968 287824
rect 66308 2176 66628 287776
rect 66968 2176 67288 287776
rect 67628 2176 67948 287776
rect 81008 2128 81328 287824
rect 81668 2176 81988 287776
rect 82328 2176 82648 287776
rect 82988 2176 83308 287776
rect 96368 2128 96688 287824
rect 97028 2176 97348 287776
rect 97688 2176 98008 287776
rect 98348 2176 98668 287776
rect 111728 2128 112048 287824
rect 112388 2176 112708 287776
rect 113048 2176 113368 287776
rect 113708 2176 114028 287776
rect 127088 2128 127408 287824
rect 127748 2176 128068 287776
rect 128408 2176 128728 287776
rect 129068 2176 129388 287776
rect 142448 2128 142768 287824
rect 143108 2176 143428 287776
rect 143768 2176 144088 287776
rect 144428 2176 144748 287776
rect 157808 2128 158128 287824
rect 158468 2176 158788 287776
rect 159128 2176 159448 287776
rect 159788 2176 160108 287776
rect 173168 2128 173488 287824
rect 173828 2176 174148 287776
rect 174488 2176 174808 287776
rect 175148 2176 175468 287776
rect 188528 2128 188848 287824
rect 189188 2176 189508 287776
rect 189848 2176 190168 287776
rect 190508 2176 190828 287776
rect 203888 2128 204208 287824
rect 204548 2176 204868 287776
rect 205208 2176 205528 287776
rect 205868 2176 206188 287776
rect 219248 2128 219568 287824
rect 219908 2176 220228 287776
rect 220568 2176 220888 287776
rect 221228 2176 221548 287776
rect 234608 2128 234928 287824
rect 235268 2176 235588 287776
rect 235928 2176 236248 287776
rect 236588 2176 236908 287776
rect 249968 2128 250288 287824
rect 250628 2176 250948 287776
rect 251288 2176 251608 287776
rect 251948 2176 252268 287776
rect 265328 2128 265648 287824
rect 265988 2176 266308 287776
rect 266648 2176 266968 287776
rect 267308 2176 267628 287776
rect 280688 2128 281008 287824
rect 281348 2176 281668 287776
rect 282008 2176 282328 287776
rect 282668 2176 282988 287776
<< obsm4 >>
rect 4659 2096 4788 287605
rect 5268 2096 5448 287605
rect 5928 2096 6108 287605
rect 6588 2096 19488 287605
rect 4659 2048 19488 2096
rect 19968 2096 20148 287605
rect 20628 2096 20808 287605
rect 21288 2096 21468 287605
rect 21948 2096 34848 287605
rect 19968 2048 34848 2096
rect 35328 2096 35508 287605
rect 35988 2096 36168 287605
rect 36648 2096 36828 287605
rect 37308 2096 50208 287605
rect 35328 2048 50208 2096
rect 50688 2096 50868 287605
rect 51348 2096 51528 287605
rect 52008 2096 52188 287605
rect 52668 2096 65568 287605
rect 50688 2048 65568 2096
rect 66048 2096 66228 287605
rect 66708 2096 66888 287605
rect 67368 2096 67548 287605
rect 68028 2096 80928 287605
rect 66048 2048 80928 2096
rect 81408 2096 81588 287605
rect 82068 2096 82248 287605
rect 82728 2096 82908 287605
rect 83388 2096 96288 287605
rect 81408 2048 96288 2096
rect 96768 2096 96948 287605
rect 97428 2096 97608 287605
rect 98088 2096 98268 287605
rect 98748 2096 111648 287605
rect 96768 2048 111648 2096
rect 112128 2096 112308 287605
rect 112788 2096 112968 287605
rect 113448 2096 113628 287605
rect 114108 2096 127008 287605
rect 112128 2048 127008 2096
rect 127488 2096 127668 287605
rect 128148 2096 128328 287605
rect 128808 2096 128988 287605
rect 129468 2096 142368 287605
rect 127488 2048 142368 2096
rect 142848 2096 143028 287605
rect 143508 2096 143688 287605
rect 144168 2096 144348 287605
rect 144828 2096 157728 287605
rect 142848 2048 157728 2096
rect 158208 2096 158388 287605
rect 158868 2096 159048 287605
rect 159528 2096 159708 287605
rect 160188 2096 173088 287605
rect 158208 2048 173088 2096
rect 173568 2096 173748 287605
rect 174228 2096 174408 287605
rect 174888 2096 175068 287605
rect 175548 2096 188448 287605
rect 173568 2048 188448 2096
rect 188928 2096 189108 287605
rect 189588 2096 189768 287605
rect 190248 2096 190428 287605
rect 190908 2096 203808 287605
rect 188928 2048 203808 2096
rect 204288 2096 204468 287605
rect 204948 2096 205128 287605
rect 205608 2096 205788 287605
rect 206268 2096 219168 287605
rect 204288 2048 219168 2096
rect 219648 2096 219828 287605
rect 220308 2096 220488 287605
rect 220968 2096 221148 287605
rect 221628 2096 234528 287605
rect 219648 2048 234528 2096
rect 235008 2096 235188 287605
rect 235668 2096 235848 287605
rect 236328 2096 236508 287605
rect 236988 2096 249888 287605
rect 235008 2048 249888 2096
rect 250368 2096 250548 287605
rect 251028 2096 251208 287605
rect 251688 2096 251868 287605
rect 252348 2096 265248 287605
rect 250368 2048 265248 2096
rect 265728 2096 265908 287605
rect 266388 2096 266568 287605
rect 267048 2096 267228 287605
rect 267708 2096 280608 287605
rect 265728 2048 280608 2096
rect 281088 2096 281268 287605
rect 281748 2096 281928 287605
rect 282408 2096 282588 287605
rect 283068 2096 289373 287605
rect 281088 2048 289373 2096
rect 4659 1259 289373 2048
<< labels >>
rlabel metal2 s 1214 289200 1270 290000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 77482 289200 77538 290000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 85118 289200 85174 290000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 92754 289200 92810 290000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 100390 289200 100446 290000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 108026 289200 108082 290000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 115662 289200 115718 290000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 123298 289200 123354 290000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 130934 289200 130990 290000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 138570 289200 138626 290000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 146206 289200 146262 290000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 8758 289200 8814 290000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 153750 289200 153806 290000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 161386 289200 161442 290000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 169022 289200 169078 290000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 176658 289200 176714 290000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 184294 289200 184350 290000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 191930 289200 191986 290000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 199566 289200 199622 290000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 207202 289200 207258 290000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 214838 289200 214894 290000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 222474 289200 222530 290000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 16394 289200 16450 290000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 230110 289200 230166 290000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 237746 289200 237802 290000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 245382 289200 245438 290000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 253018 289200 253074 290000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 260654 289200 260710 290000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 268290 289200 268346 290000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 275926 289200 275982 290000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 283562 289200 283618 290000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 24030 289200 24086 290000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 31666 289200 31722 290000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 39302 289200 39358 290000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 46938 289200 46994 290000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 54574 289200 54630 290000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 62210 289200 62266 290000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 69846 289200 69902 290000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3698 289200 3754 290000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 80058 289200 80114 290000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 87694 289200 87750 290000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 95330 289200 95386 290000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 102874 289200 102930 290000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 110510 289200 110566 290000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 118146 289200 118202 290000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 125782 289200 125838 290000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 133418 289200 133474 290000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 141054 289200 141110 290000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 148690 289200 148746 290000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 11334 289200 11390 290000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 156326 289200 156382 290000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 163962 289200 164018 290000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 171598 289200 171654 290000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 179234 289200 179290 290000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 186870 289200 186926 290000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 194506 289200 194562 290000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 202142 289200 202198 290000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 209778 289200 209834 290000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 217414 289200 217470 290000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 225050 289200 225106 290000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 18970 289200 19026 290000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 232686 289200 232742 290000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 240322 289200 240378 290000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 247866 289200 247922 290000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 255502 289200 255558 290000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 263138 289200 263194 290000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 270774 289200 270830 290000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 278410 289200 278466 290000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 286046 289200 286102 290000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 26606 289200 26662 290000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 34242 289200 34298 290000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 41878 289200 41934 290000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 49514 289200 49570 290000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 57150 289200 57206 290000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 64786 289200 64842 290000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 72422 289200 72478 290000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 6274 289200 6330 290000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 82542 289200 82598 290000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 90178 289200 90234 290000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 97814 289200 97870 290000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 105450 289200 105506 290000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 113086 289200 113142 290000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 120722 289200 120778 290000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 128358 289200 128414 290000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 135994 289200 136050 290000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 143630 289200 143686 290000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 151266 289200 151322 290000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 13910 289200 13966 290000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 158902 289200 158958 290000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 166538 289200 166594 290000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 174174 289200 174230 290000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 181810 289200 181866 290000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 189446 289200 189502 290000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 196990 289200 197046 290000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 204626 289200 204682 290000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 212262 289200 212318 290000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 219898 289200 219954 290000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 227534 289200 227590 290000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 21546 289200 21602 290000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 235170 289200 235226 290000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 242806 289200 242862 290000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 250442 289200 250498 290000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 258078 289200 258134 290000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 265714 289200 265770 290000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 273350 289200 273406 290000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 280986 289200 281042 290000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 288622 289200 288678 290000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 29182 289200 29238 290000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 36818 289200 36874 290000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 44454 289200 44510 290000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 51998 289200 52054 290000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 59634 289200 59690 290000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 67270 289200 67326 290000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 74906 289200 74962 290000 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 289200 217472 290000 217592 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 0 144984 800 145104 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 289634 0 289690 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 240046 0 240102 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 241794 0 241850 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 243542 0 243598 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 245382 0 245438 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 247130 0 247186 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 248878 0 248934 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 250626 0 250682 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 252466 0 252522 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 254214 0 254270 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 255962 0 256018 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 257710 0 257766 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 259550 0 259606 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 261298 0 261354 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 263046 0 263102 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 264794 0 264850 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 266634 0 266690 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 268382 0 268438 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 270130 0 270186 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 271878 0 271934 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 273718 0 273774 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 275466 0 275522 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 277214 0 277270 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 279054 0 279110 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 280802 0 280858 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 282550 0 282606 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 284298 0 284354 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 286138 0 286194 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 287886 0 287942 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 128450 0 128506 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 131946 0 132002 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 133694 0 133750 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 139030 0 139086 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 140778 0 140834 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 144366 0 144422 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 146114 0 146170 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 147862 0 147918 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 149702 0 149758 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 151450 0 151506 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 156786 0 156842 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 158534 0 158590 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 160282 0 160338 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 162030 0 162086 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 163870 0 163926 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 165618 0 165674 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 167366 0 167422 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 172702 0 172758 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 174450 0 174506 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 176290 0 176346 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 178038 0 178094 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 179786 0 179842 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 181534 0 181590 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 183374 0 183430 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 185122 0 185178 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 186870 0 186926 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 188618 0 188674 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 190458 0 190514 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 192206 0 192262 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 193954 0 194010 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 195702 0 195758 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 197542 0 197598 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 199290 0 199346 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 201038 0 201094 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 202786 0 202842 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 204626 0 204682 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 206374 0 206430 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 208122 0 208178 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 209870 0 209926 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 211710 0 211766 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 213458 0 213514 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 215206 0 215262 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 216954 0 217010 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 218794 0 218850 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 220542 0 220598 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 222290 0 222346 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 224130 0 224186 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 225878 0 225934 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 227626 0 227682 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 229374 0 229430 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 231214 0 231270 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 232962 0 233018 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 234710 0 234766 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 236458 0 236514 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 238298 0 238354 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 240598 0 240654 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 242438 0 242494 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 244186 0 244242 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 245934 0 245990 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 247682 0 247738 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 249522 0 249578 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 251270 0 251326 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 253018 0 253074 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 254766 0 254822 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 256606 0 256662 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 258354 0 258410 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 260102 0 260158 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 261850 0 261906 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 263690 0 263746 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 265438 0 265494 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 267186 0 267242 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 268934 0 268990 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 270774 0 270830 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 272522 0 272578 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 274270 0 274326 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 82910 0 82966 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 276018 0 276074 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 277858 0 277914 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 279606 0 279662 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 281354 0 281410 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 283102 0 283158 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 284942 0 284998 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 286690 0 286746 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 288438 0 288494 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 89994 0 90050 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 91834 0 91890 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 93582 0 93638 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 97078 0 97134 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 100666 0 100722 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 102414 0 102470 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 104162 0 104218 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 106002 0 106058 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 107750 0 107806 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 111246 0 111302 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 113086 0 113142 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 114834 0 114890 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 118330 0 118386 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 120170 0 120226 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 125414 0 125470 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 127254 0 127310 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 132498 0 132554 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 134338 0 134394 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 136086 0 136142 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 137834 0 137890 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 139674 0 139730 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 141422 0 141478 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 143170 0 143226 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 146758 0 146814 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 148506 0 148562 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 150254 0 150310 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 152002 0 152058 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 153842 0 153898 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 155590 0 155646 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 157338 0 157394 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 159086 0 159142 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 160926 0 160982 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 162674 0 162730 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 164422 0 164478 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 166170 0 166226 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 168010 0 168066 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 72330 0 72386 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 169758 0 169814 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 171506 0 171562 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 173254 0 173310 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 175094 0 175150 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 176842 0 176898 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 178590 0 178646 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 180338 0 180394 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 182178 0 182234 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 183926 0 183982 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 185674 0 185730 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 187422 0 187478 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 189262 0 189318 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 191010 0 191066 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 192758 0 192814 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 194598 0 194654 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 196346 0 196402 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 198094 0 198150 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 199842 0 199898 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 201682 0 201738 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 203430 0 203486 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 75826 0 75882 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 205178 0 205234 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 206926 0 206982 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 208766 0 208822 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 210514 0 210570 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 212262 0 212318 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 214010 0 214066 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 215850 0 215906 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 217598 0 217654 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 219346 0 219402 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 221094 0 221150 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 222934 0 222990 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 224682 0 224738 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 226430 0 226486 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 228178 0 228234 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 230018 0 230074 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 231766 0 231822 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 233514 0 233570 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 235262 0 235318 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 237102 0 237158 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 238850 0 238906 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 64050 0 64106 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 241242 0 241298 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 242990 0 243046 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 244738 0 244794 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 246486 0 246542 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 248326 0 248382 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 250074 0 250130 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 251822 0 251878 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 253570 0 253626 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 255410 0 255466 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 257158 0 257214 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 258906 0 258962 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 260746 0 260802 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 262494 0 262550 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 264242 0 264298 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 265990 0 266046 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 267830 0 267886 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 269578 0 269634 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 271326 0 271382 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 273074 0 273130 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 274914 0 274970 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 276662 0 276718 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 278410 0 278466 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 280158 0 280214 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 281998 0 282054 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 283746 0 283802 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 285494 0 285550 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 287242 0 287298 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 289082 0 289138 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 106554 0 106610 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 122470 0 122526 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 126058 0 126114 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 129554 0 129610 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 140226 0 140282 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 141974 0 142030 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 147310 0 147366 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 150806 0 150862 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 152646 0 152702 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 156142 0 156198 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 161478 0 161534 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 163226 0 163282 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 166814 0 166870 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 168562 0 168618 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 170310 0 170366 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 172150 0 172206 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 173898 0 173954 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 175646 0 175702 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 177394 0 177450 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 179234 0 179290 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 182730 0 182786 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 184478 0 184534 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 186318 0 186374 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 188066 0 188122 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 189814 0 189870 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 191562 0 191618 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 193402 0 193458 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 195150 0 195206 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 196898 0 196954 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 198646 0 198702 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 200486 0 200542 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 202234 0 202290 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 203982 0 204038 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 205822 0 205878 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 207570 0 207626 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 209318 0 209374 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 211066 0 211122 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 212906 0 212962 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 214654 0 214710 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 216402 0 216458 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 218150 0 218206 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 219990 0 220046 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 221738 0 221794 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 223486 0 223542 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 225234 0 225290 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 227074 0 227130 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 228822 0 228878 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 230570 0 230626 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 232318 0 232374 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 234158 0 234214 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 235906 0 235962 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 237654 0 237710 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 239402 0 239458 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal3 s 289200 72496 290000 72616 6 user_clk
port 502 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 503 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 504 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_ack_o
port 505 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 wbs_adr_i[0]
port 506 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_adr_i[10]
port 507 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_adr_i[11]
port 508 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wbs_adr_i[12]
port 509 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_adr_i[13]
port 510 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wbs_adr_i[14]
port 511 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_adr_i[15]
port 512 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 wbs_adr_i[16]
port 513 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 wbs_adr_i[17]
port 514 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_adr_i[18]
port 515 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 wbs_adr_i[19]
port 516 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_adr_i[1]
port 517 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 wbs_adr_i[20]
port 518 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 wbs_adr_i[21]
port 519 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 wbs_adr_i[22]
port 520 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 wbs_adr_i[23]
port 521 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 wbs_adr_i[24]
port 522 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 wbs_adr_i[25]
port 523 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 wbs_adr_i[26]
port 524 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 wbs_adr_i[27]
port 525 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 wbs_adr_i[28]
port 526 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 wbs_adr_i[29]
port 527 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[2]
port 528 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 wbs_adr_i[30]
port 529 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 wbs_adr_i[31]
port 530 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_adr_i[3]
port 531 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_adr_i[4]
port 532 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_adr_i[5]
port 533 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[6]
port 534 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[7]
port 535 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[8]
port 536 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_adr_i[9]
port 537 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_cyc_i
port 538 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_i[0]
port 539 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_dat_i[10]
port 540 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_i[11]
port 541 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_i[12]
port 542 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_dat_i[13]
port 543 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_i[14]
port 544 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_i[15]
port 545 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 wbs_dat_i[16]
port 546 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_i[17]
port 547 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_i[18]
port 548 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 wbs_dat_i[19]
port 549 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_i[1]
port 550 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 wbs_dat_i[20]
port 551 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 wbs_dat_i[21]
port 552 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wbs_dat_i[22]
port 553 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 wbs_dat_i[23]
port 554 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 wbs_dat_i[24]
port 555 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 wbs_dat_i[25]
port 556 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 wbs_dat_i[26]
port 557 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 wbs_dat_i[27]
port 558 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 wbs_dat_i[28]
port 559 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 wbs_dat_i[29]
port 560 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_dat_i[2]
port 561 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 wbs_dat_i[30]
port 562 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 wbs_dat_i[31]
port 563 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[3]
port 564 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[4]
port 565 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_i[5]
port 566 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_i[6]
port 567 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_dat_i[7]
port 568 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_i[8]
port 569 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_dat_i[9]
port 570 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_o[0]
port 571 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_o[10]
port 572 nsew signal output
rlabel metal2 s 26790 0 26846 800 6 wbs_dat_o[11]
port 573 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_o[12]
port 574 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_o[13]
port 575 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_o[14]
port 576 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_o[15]
port 577 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 wbs_dat_o[16]
port 578 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_o[17]
port 579 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 wbs_dat_o[18]
port 580 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 wbs_dat_o[19]
port 581 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[1]
port 582 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_o[20]
port 583 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 wbs_dat_o[21]
port 584 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 wbs_dat_o[22]
port 585 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 wbs_dat_o[23]
port 586 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 wbs_dat_o[24]
port 587 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 wbs_dat_o[25]
port 588 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 wbs_dat_o[26]
port 589 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 wbs_dat_o[27]
port 590 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 wbs_dat_o[28]
port 591 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 wbs_dat_o[29]
port 592 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_o[2]
port 593 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 wbs_dat_o[30]
port 594 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 wbs_dat_o[31]
port 595 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_o[3]
port 596 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_o[4]
port 597 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_o[5]
port 598 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 wbs_dat_o[6]
port 599 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_o[7]
port 600 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_o[8]
port 601 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_o[9]
port 602 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wbs_sel_i[0]
port 603 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_sel_i[1]
port 604 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_sel_i[2]
port 605 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_sel_i[3]
port 606 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_stb_i
port 607 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_we_i
port 608 nsew signal input
rlabel metal4 s 280688 2128 281008 287824 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 287824 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 287824 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 287824 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 287824 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 287824 6 vccd1
port 614 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 287824 6 vccd1
port 615 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 287824 6 vccd1
port 616 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 287824 6 vccd1
port 617 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 287824 6 vccd1
port 618 nsew power bidirectional
rlabel metal4 s 265328 2128 265648 287824 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 287824 6 vssd1
port 620 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 287824 6 vssd1
port 621 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 287824 6 vssd1
port 622 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 287824 6 vssd1
port 623 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 287824 6 vssd1
port 624 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 287824 6 vssd1
port 625 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 287824 6 vssd1
port 626 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 287824 6 vssd1
port 627 nsew ground bidirectional
rlabel metal4 s 281348 2176 281668 287776 6 vccd2
port 628 nsew power bidirectional
rlabel metal4 s 250628 2176 250948 287776 6 vccd2
port 629 nsew power bidirectional
rlabel metal4 s 219908 2176 220228 287776 6 vccd2
port 630 nsew power bidirectional
rlabel metal4 s 189188 2176 189508 287776 6 vccd2
port 631 nsew power bidirectional
rlabel metal4 s 158468 2176 158788 287776 6 vccd2
port 632 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 287776 6 vccd2
port 633 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 287776 6 vccd2
port 634 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 287776 6 vccd2
port 635 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 287776 6 vccd2
port 636 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 287776 6 vccd2
port 637 nsew power bidirectional
rlabel metal4 s 265988 2176 266308 287776 6 vssd2
port 638 nsew ground bidirectional
rlabel metal4 s 235268 2176 235588 287776 6 vssd2
port 639 nsew ground bidirectional
rlabel metal4 s 204548 2176 204868 287776 6 vssd2
port 640 nsew ground bidirectional
rlabel metal4 s 173828 2176 174148 287776 6 vssd2
port 641 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 287776 6 vssd2
port 642 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 287776 6 vssd2
port 643 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 287776 6 vssd2
port 644 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 287776 6 vssd2
port 645 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 287776 6 vssd2
port 646 nsew ground bidirectional
rlabel metal4 s 282008 2176 282328 287776 6 vdda1
port 647 nsew power bidirectional
rlabel metal4 s 251288 2176 251608 287776 6 vdda1
port 648 nsew power bidirectional
rlabel metal4 s 220568 2176 220888 287776 6 vdda1
port 649 nsew power bidirectional
rlabel metal4 s 189848 2176 190168 287776 6 vdda1
port 650 nsew power bidirectional
rlabel metal4 s 159128 2176 159448 287776 6 vdda1
port 651 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 287776 6 vdda1
port 652 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 287776 6 vdda1
port 653 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 287776 6 vdda1
port 654 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 287776 6 vdda1
port 655 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 287776 6 vdda1
port 656 nsew power bidirectional
rlabel metal4 s 266648 2176 266968 287776 6 vssa1
port 657 nsew ground bidirectional
rlabel metal4 s 235928 2176 236248 287776 6 vssa1
port 658 nsew ground bidirectional
rlabel metal4 s 205208 2176 205528 287776 6 vssa1
port 659 nsew ground bidirectional
rlabel metal4 s 174488 2176 174808 287776 6 vssa1
port 660 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 287776 6 vssa1
port 661 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 287776 6 vssa1
port 662 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 287776 6 vssa1
port 663 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 287776 6 vssa1
port 664 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 287776 6 vssa1
port 665 nsew ground bidirectional
rlabel metal4 s 282668 2176 282988 287776 6 vdda2
port 666 nsew power bidirectional
rlabel metal4 s 251948 2176 252268 287776 6 vdda2
port 667 nsew power bidirectional
rlabel metal4 s 221228 2176 221548 287776 6 vdda2
port 668 nsew power bidirectional
rlabel metal4 s 190508 2176 190828 287776 6 vdda2
port 669 nsew power bidirectional
rlabel metal4 s 159788 2176 160108 287776 6 vdda2
port 670 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 287776 6 vdda2
port 671 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 287776 6 vdda2
port 672 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 287776 6 vdda2
port 673 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 287776 6 vdda2
port 674 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 287776 6 vdda2
port 675 nsew power bidirectional
rlabel metal4 s 267308 2176 267628 287776 6 vssa2
port 676 nsew ground bidirectional
rlabel metal4 s 236588 2176 236908 287776 6 vssa2
port 677 nsew ground bidirectional
rlabel metal4 s 205868 2176 206188 287776 6 vssa2
port 678 nsew ground bidirectional
rlabel metal4 s 175148 2176 175468 287776 6 vssa2
port 679 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 287776 6 vssa2
port 680 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 287776 6 vssa2
port 681 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 287776 6 vssa2
port 682 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 287776 6 vssa2
port 683 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 287776 6 vssa2
port 684 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 290000 290000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj.gds
string GDS_END 269490638
string GDS_START 843676
<< end >>

