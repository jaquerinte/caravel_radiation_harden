VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 1490.000 BY 1490.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 1486.000 6.350 1490.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 1486.000 391.370 1490.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 1486.000 430.010 1490.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 1486.000 468.650 1490.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 1486.000 506.830 1490.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 1486.000 545.470 1490.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 1486.000 584.110 1490.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 1486.000 622.750 1490.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 1486.000 661.390 1490.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 1486.000 699.570 1490.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 1486.000 738.210 1490.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 1486.000 44.530 1490.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 1486.000 776.850 1490.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 1486.000 815.490 1490.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 1486.000 853.670 1490.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 1486.000 892.310 1490.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.670 1486.000 930.950 1490.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 1486.000 969.590 1490.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.490 1486.000 1007.770 1490.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.130 1486.000 1046.410 1490.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.770 1486.000 1085.050 1490.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.410 1486.000 1123.690 1490.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 1486.000 83.170 1490.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.050 1486.000 1162.330 1490.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1200.230 1486.000 1200.510 1490.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.870 1486.000 1239.150 1490.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.510 1486.000 1277.790 1490.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.150 1486.000 1316.430 1490.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1354.330 1486.000 1354.610 1490.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.970 1486.000 1393.250 1490.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.610 1486.000 1431.890 1490.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 1486.000 121.810 1490.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 1486.000 160.450 1490.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 1486.000 198.630 1490.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 1486.000 237.270 1490.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 1486.000 275.910 1490.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 1486.000 314.550 1490.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 1486.000 352.730 1490.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 1486.000 18.770 1490.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 1486.000 404.250 1490.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 1486.000 442.890 1490.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 1486.000 481.530 1490.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 1486.000 519.710 1490.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 1486.000 558.350 1490.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.710 1486.000 596.990 1490.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 1486.000 635.630 1490.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 1486.000 673.810 1490.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 1486.000 712.450 1490.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 1486.000 751.090 1490.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 1486.000 57.410 1490.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 1486.000 789.730 1490.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 1486.000 828.370 1490.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 1486.000 866.550 1490.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 1486.000 905.190 1490.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 1486.000 943.830 1490.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 1486.000 982.470 1490.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.370 1486.000 1020.650 1490.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.010 1486.000 1059.290 1490.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.650 1486.000 1097.930 1490.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.290 1486.000 1136.570 1490.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 1486.000 96.050 1490.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.470 1486.000 1174.750 1490.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1213.110 1486.000 1213.390 1490.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.750 1486.000 1252.030 1490.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1290.390 1486.000 1290.670 1490.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.030 1486.000 1329.310 1490.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.210 1486.000 1367.490 1490.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.850 1486.000 1406.130 1490.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.490 1486.000 1444.770 1490.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 1486.000 134.690 1490.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 1486.000 172.870 1490.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 1486.000 211.510 1490.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 1486.000 250.150 1490.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 1486.000 288.790 1490.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 1486.000 327.430 1490.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 1486.000 365.610 1490.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 1486.000 31.650 1490.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 1486.000 417.130 1490.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 1486.000 455.770 1490.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 1486.000 494.410 1490.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 1486.000 532.590 1490.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 1486.000 571.230 1490.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 1486.000 609.870 1490.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.230 1486.000 648.510 1490.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 1486.000 686.690 1490.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 1486.000 725.330 1490.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 1486.000 763.970 1490.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 1486.000 70.290 1490.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 1486.000 802.610 1490.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 1486.000 840.790 1490.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 1486.000 879.430 1490.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 1486.000 918.070 1490.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 1486.000 956.710 1490.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 1486.000 995.350 1490.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.250 1486.000 1033.530 1490.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.890 1486.000 1072.170 1490.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.530 1486.000 1110.810 1490.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.170 1486.000 1149.450 1490.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 1486.000 108.930 1490.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.350 1486.000 1187.630 1490.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.990 1486.000 1226.270 1490.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.630 1486.000 1264.910 1490.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.270 1486.000 1303.550 1490.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1341.450 1486.000 1341.730 1490.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.090 1486.000 1380.370 1490.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.730 1486.000 1419.010 1490.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1457.370 1486.000 1457.650 1490.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 1486.000 147.570 1490.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 1486.000 185.750 1490.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 1486.000 224.390 1490.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 1486.000 263.030 1490.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 1486.000 301.670 1490.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 1486.000 339.850 1490.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 1486.000 378.490 1490.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 0.000 744.640 4.000 745.240 ;
=======
      LAYER met2 ;
        RECT 895.250 0.000 895.530 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1470.250 1486.000 1470.530 1490.000 ;
=======
        RECT 897.090 0.000 897.370 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1483.130 1486.000 1483.410 1490.000 ;
=======
        RECT 898.930 0.000 899.210 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 323.010 0.000 323.290 4.000 ;
=======
        RECT 193.750 0.000 194.030 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1233.350 0.000 1233.630 4.000 ;
=======
        RECT 741.610 0.000 741.890 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1242.550 0.000 1242.830 4.000 ;
=======
        RECT 747.130 0.000 747.410 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1251.290 0.000 1251.570 4.000 ;
=======
        RECT 752.650 0.000 752.930 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1260.490 0.000 1260.770 4.000 ;
=======
        RECT 758.170 0.000 758.450 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1269.690 0.000 1269.970 4.000 ;
=======
        RECT 763.690 0.000 763.970 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1278.890 0.000 1279.170 4.000 ;
=======
        RECT 769.210 0.000 769.490 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1288.090 0.000 1288.370 4.000 ;
=======
        RECT 774.730 0.000 775.010 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1296.830 0.000 1297.110 4.000 ;
=======
        RECT 780.250 0.000 780.530 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1306.030 0.000 1306.310 4.000 ;
=======
        RECT 785.310 0.000 785.590 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1315.230 0.000 1315.510 4.000 ;
=======
        RECT 790.830 0.000 791.110 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 414.090 0.000 414.370 4.000 ;
=======
        RECT 248.490 0.000 248.770 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1324.430 0.000 1324.710 4.000 ;
=======
        RECT 796.350 0.000 796.630 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1333.170 0.000 1333.450 4.000 ;
=======
        RECT 801.870 0.000 802.150 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1342.370 0.000 1342.650 4.000 ;
=======
        RECT 807.390 0.000 807.670 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1351.570 0.000 1351.850 4.000 ;
=======
        RECT 812.910 0.000 813.190 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1360.770 0.000 1361.050 4.000 ;
=======
        RECT 818.430 0.000 818.710 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1369.970 0.000 1370.250 4.000 ;
=======
        RECT 823.950 0.000 824.230 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1378.710 0.000 1378.990 4.000 ;
=======
        RECT 829.470 0.000 829.750 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1387.910 0.000 1388.190 4.000 ;
=======
        RECT 834.990 0.000 835.270 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1397.110 0.000 1397.390 4.000 ;
=======
        RECT 840.510 0.000 840.790 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1406.310 0.000 1406.590 4.000 ;
=======
        RECT 845.570 0.000 845.850 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 422.830 0.000 423.110 4.000 ;
=======
        RECT 254.010 0.000 254.290 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1415.510 0.000 1415.790 4.000 ;
=======
        RECT 851.090 0.000 851.370 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1424.250 0.000 1424.530 4.000 ;
=======
        RECT 856.610 0.000 856.890 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1433.450 0.000 1433.730 4.000 ;
=======
        RECT 862.130 0.000 862.410 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1442.650 0.000 1442.930 4.000 ;
=======
        RECT 867.650 0.000 867.930 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1451.850 0.000 1452.130 4.000 ;
=======
        RECT 873.170 0.000 873.450 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1461.050 0.000 1461.330 4.000 ;
=======
        RECT 878.690 0.000 878.970 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1469.790 0.000 1470.070 4.000 ;
=======
        RECT 884.210 0.000 884.490 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1478.990 0.000 1479.270 4.000 ;
=======
        RECT 889.730 0.000 890.010 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 432.030 0.000 432.310 4.000 ;
=======
        RECT 259.530 0.000 259.810 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 441.230 0.000 441.510 4.000 ;
=======
        RECT 265.050 0.000 265.330 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 450.430 0.000 450.710 4.000 ;
=======
        RECT 270.570 0.000 270.850 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 459.630 0.000 459.910 4.000 ;
=======
        RECT 276.090 0.000 276.370 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 468.370 0.000 468.650 4.000 ;
=======
        RECT 281.610 0.000 281.890 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 477.570 0.000 477.850 4.000 ;
=======
        RECT 287.130 0.000 287.410 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 486.770 0.000 487.050 4.000 ;
=======
        RECT 292.650 0.000 292.930 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 495.970 0.000 496.250 4.000 ;
=======
        RECT 298.170 0.000 298.450 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 332.210 0.000 332.490 4.000 ;
=======
        RECT 199.270 0.000 199.550 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 505.170 0.000 505.450 4.000 ;
=======
        RECT 303.230 0.000 303.510 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 513.910 0.000 514.190 4.000 ;
=======
        RECT 308.750 0.000 309.030 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 523.110 0.000 523.390 4.000 ;
=======
        RECT 314.270 0.000 314.550 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 532.310 0.000 532.590 4.000 ;
=======
        RECT 319.790 0.000 320.070 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 541.510 0.000 541.790 4.000 ;
=======
        RECT 325.310 0.000 325.590 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 550.710 0.000 550.990 4.000 ;
=======
        RECT 330.830 0.000 331.110 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 559.450 0.000 559.730 4.000 ;
=======
        RECT 336.350 0.000 336.630 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 568.650 0.000 568.930 4.000 ;
=======
        RECT 341.870 0.000 342.150 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 577.850 0.000 578.130 4.000 ;
=======
        RECT 347.390 0.000 347.670 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 587.050 0.000 587.330 4.000 ;
=======
        RECT 352.910 0.000 353.190 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 340.950 0.000 341.230 4.000 ;
=======
        RECT 204.790 0.000 205.070 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 595.790 0.000 596.070 4.000 ;
=======
        RECT 358.430 0.000 358.710 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 604.990 0.000 605.270 4.000 ;
=======
        RECT 363.490 0.000 363.770 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 614.190 0.000 614.470 4.000 ;
=======
        RECT 369.010 0.000 369.290 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 623.390 0.000 623.670 4.000 ;
=======
        RECT 374.530 0.000 374.810 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 632.590 0.000 632.870 4.000 ;
=======
        RECT 380.050 0.000 380.330 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 641.330 0.000 641.610 4.000 ;
=======
        RECT 385.570 0.000 385.850 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 650.530 0.000 650.810 4.000 ;
=======
        RECT 391.090 0.000 391.370 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 659.730 0.000 660.010 4.000 ;
=======
        RECT 396.610 0.000 396.890 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 668.930 0.000 669.210 4.000 ;
=======
        RECT 402.130 0.000 402.410 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 678.130 0.000 678.410 4.000 ;
=======
        RECT 407.650 0.000 407.930 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 350.150 0.000 350.430 4.000 ;
=======
        RECT 210.310 0.000 210.590 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 686.870 0.000 687.150 4.000 ;
=======
        RECT 413.170 0.000 413.450 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 696.070 0.000 696.350 4.000 ;
=======
        RECT 418.690 0.000 418.970 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 705.270 0.000 705.550 4.000 ;
=======
        RECT 423.750 0.000 424.030 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 714.470 0.000 714.750 4.000 ;
=======
        RECT 429.270 0.000 429.550 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 723.670 0.000 723.950 4.000 ;
=======
        RECT 434.790 0.000 435.070 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 732.410 0.000 732.690 4.000 ;
=======
        RECT 440.310 0.000 440.590 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 741.610 0.000 741.890 4.000 ;
=======
        RECT 445.830 0.000 446.110 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 750.810 0.000 751.090 4.000 ;
=======
        RECT 451.350 0.000 451.630 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 760.010 0.000 760.290 4.000 ;
=======
        RECT 456.870 0.000 457.150 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 768.750 0.000 769.030 4.000 ;
=======
        RECT 462.390 0.000 462.670 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 359.350 0.000 359.630 4.000 ;
=======
        RECT 215.830 0.000 216.110 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 777.950 0.000 778.230 4.000 ;
=======
        RECT 467.910 0.000 468.190 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 787.150 0.000 787.430 4.000 ;
=======
        RECT 473.430 0.000 473.710 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 796.350 0.000 796.630 4.000 ;
=======
        RECT 478.950 0.000 479.230 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 805.550 0.000 805.830 4.000 ;
=======
        RECT 484.010 0.000 484.290 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 814.290 0.000 814.570 4.000 ;
=======
        RECT 489.530 0.000 489.810 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 823.490 0.000 823.770 4.000 ;
=======
        RECT 495.050 0.000 495.330 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 832.690 0.000 832.970 4.000 ;
=======
        RECT 500.570 0.000 500.850 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 841.890 0.000 842.170 4.000 ;
=======
        RECT 506.090 0.000 506.370 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 851.090 0.000 851.370 4.000 ;
=======
        RECT 511.610 0.000 511.890 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 859.830 0.000 860.110 4.000 ;
=======
        RECT 517.130 0.000 517.410 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 368.550 0.000 368.830 4.000 ;
=======
        RECT 221.350 0.000 221.630 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 869.030 0.000 869.310 4.000 ;
=======
        RECT 522.650 0.000 522.930 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 878.230 0.000 878.510 4.000 ;
=======
        RECT 528.170 0.000 528.450 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 887.430 0.000 887.710 4.000 ;
=======
        RECT 533.690 0.000 533.970 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 896.630 0.000 896.910 4.000 ;
=======
        RECT 539.210 0.000 539.490 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 905.370 0.000 905.650 4.000 ;
=======
        RECT 544.270 0.000 544.550 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 914.570 0.000 914.850 4.000 ;
=======
        RECT 549.790 0.000 550.070 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 923.770 0.000 924.050 4.000 ;
=======
        RECT 555.310 0.000 555.590 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 932.970 0.000 933.250 4.000 ;
=======
        RECT 560.830 0.000 561.110 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 941.710 0.000 941.990 4.000 ;
=======
        RECT 566.350 0.000 566.630 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 950.910 0.000 951.190 4.000 ;
=======
        RECT 571.870 0.000 572.150 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 377.290 0.000 377.570 4.000 ;
=======
        RECT 226.870 0.000 227.150 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 960.110 0.000 960.390 4.000 ;
=======
        RECT 577.390 0.000 577.670 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 969.310 0.000 969.590 4.000 ;
=======
        RECT 582.910 0.000 583.190 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 978.510 0.000 978.790 4.000 ;
=======
        RECT 588.430 0.000 588.710 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 987.250 0.000 987.530 4.000 ;
=======
        RECT 593.950 0.000 594.230 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 996.450 0.000 996.730 4.000 ;
=======
        RECT 599.470 0.000 599.750 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1005.650 0.000 1005.930 4.000 ;
=======
        RECT 604.530 0.000 604.810 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1014.850 0.000 1015.130 4.000 ;
=======
        RECT 610.050 0.000 610.330 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1024.050 0.000 1024.330 4.000 ;
=======
        RECT 615.570 0.000 615.850 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1032.790 0.000 1033.070 4.000 ;
=======
        RECT 621.090 0.000 621.370 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1041.990 0.000 1042.270 4.000 ;
=======
        RECT 626.610 0.000 626.890 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 386.490 0.000 386.770 4.000 ;
=======
        RECT 232.390 0.000 232.670 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1051.190 0.000 1051.470 4.000 ;
=======
        RECT 632.130 0.000 632.410 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1060.390 0.000 1060.670 4.000 ;
=======
        RECT 637.650 0.000 637.930 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1069.590 0.000 1069.870 4.000 ;
=======
        RECT 643.170 0.000 643.450 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1078.330 0.000 1078.610 4.000 ;
=======
        RECT 648.690 0.000 648.970 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1087.530 0.000 1087.810 4.000 ;
=======
        RECT 654.210 0.000 654.490 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1096.730 0.000 1097.010 4.000 ;
=======
        RECT 659.730 0.000 660.010 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1105.930 0.000 1106.210 4.000 ;
=======
        RECT 664.790 0.000 665.070 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1115.130 0.000 1115.410 4.000 ;
=======
        RECT 670.310 0.000 670.590 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1123.870 0.000 1124.150 4.000 ;
=======
        RECT 675.830 0.000 676.110 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1133.070 0.000 1133.350 4.000 ;
=======
        RECT 681.350 0.000 681.630 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 395.690 0.000 395.970 4.000 ;
=======
        RECT 237.910 0.000 238.190 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1142.270 0.000 1142.550 4.000 ;
=======
        RECT 686.870 0.000 687.150 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1151.470 0.000 1151.750 4.000 ;
=======
        RECT 692.390 0.000 692.670 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1160.210 0.000 1160.490 4.000 ;
=======
        RECT 697.910 0.000 698.190 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1169.410 0.000 1169.690 4.000 ;
=======
        RECT 703.430 0.000 703.710 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1178.610 0.000 1178.890 4.000 ;
=======
        RECT 708.950 0.000 709.230 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1187.810 0.000 1188.090 4.000 ;
=======
        RECT 714.470 0.000 714.750 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1197.010 0.000 1197.290 4.000 ;
=======
        RECT 719.990 0.000 720.270 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1205.750 0.000 1206.030 4.000 ;
=======
        RECT 725.050 0.000 725.330 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1214.950 0.000 1215.230 4.000 ;
=======
        RECT 730.570 0.000 730.850 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1224.150 0.000 1224.430 4.000 ;
=======
        RECT 736.090 0.000 736.370 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 404.890 0.000 405.170 4.000 ;
=======
        RECT 242.970 0.000 243.250 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 325.770 0.000 326.050 4.000 ;
=======
        RECT 195.590 0.000 195.870 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1236.110 0.000 1236.390 4.000 ;
=======
        RECT 743.450 0.000 743.730 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1245.310 0.000 1245.590 4.000 ;
=======
        RECT 748.970 0.000 749.250 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1254.510 0.000 1254.790 4.000 ;
=======
        RECT 754.490 0.000 754.770 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1263.710 0.000 1263.990 4.000 ;
=======
        RECT 760.010 0.000 760.290 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1272.910 0.000 1273.190 4.000 ;
=======
        RECT 765.530 0.000 765.810 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1281.650 0.000 1281.930 4.000 ;
=======
        RECT 771.050 0.000 771.330 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1290.850 0.000 1291.130 4.000 ;
=======
        RECT 776.570 0.000 776.850 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1300.050 0.000 1300.330 4.000 ;
=======
        RECT 781.630 0.000 781.910 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1309.250 0.000 1309.530 4.000 ;
=======
        RECT 787.150 0.000 787.430 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1317.990 0.000 1318.270 4.000 ;
=======
        RECT 792.670 0.000 792.950 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 416.850 0.000 417.130 4.000 ;
=======
        RECT 250.330 0.000 250.610 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1327.190 0.000 1327.470 4.000 ;
=======
        RECT 798.190 0.000 798.470 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1336.390 0.000 1336.670 4.000 ;
=======
        RECT 803.710 0.000 803.990 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1345.590 0.000 1345.870 4.000 ;
=======
        RECT 809.230 0.000 809.510 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1354.790 0.000 1355.070 4.000 ;
=======
        RECT 814.750 0.000 815.030 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1363.530 0.000 1363.810 4.000 ;
=======
        RECT 820.270 0.000 820.550 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1372.730 0.000 1373.010 4.000 ;
=======
        RECT 825.790 0.000 826.070 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1381.930 0.000 1382.210 4.000 ;
=======
        RECT 831.310 0.000 831.590 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1391.130 0.000 1391.410 4.000 ;
=======
        RECT 836.830 0.000 837.110 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1400.330 0.000 1400.610 4.000 ;
=======
        RECT 841.890 0.000 842.170 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1409.070 0.000 1409.350 4.000 ;
=======
        RECT 847.410 0.000 847.690 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 426.050 0.000 426.330 4.000 ;
=======
        RECT 255.850 0.000 256.130 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1418.270 0.000 1418.550 4.000 ;
=======
        RECT 852.930 0.000 853.210 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1427.470 0.000 1427.750 4.000 ;
=======
        RECT 858.450 0.000 858.730 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1436.670 0.000 1436.950 4.000 ;
=======
        RECT 863.970 0.000 864.250 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1445.870 0.000 1446.150 4.000 ;
=======
        RECT 869.490 0.000 869.770 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1454.610 0.000 1454.890 4.000 ;
=======
        RECT 875.010 0.000 875.290 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1463.810 0.000 1464.090 4.000 ;
=======
        RECT 880.530 0.000 880.810 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1473.010 0.000 1473.290 4.000 ;
=======
        RECT 886.050 0.000 886.330 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1482.210 0.000 1482.490 4.000 ;
=======
        RECT 891.570 0.000 891.850 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 435.250 0.000 435.530 4.000 ;
=======
        RECT 261.370 0.000 261.650 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 444.450 0.000 444.730 4.000 ;
=======
        RECT 266.890 0.000 267.170 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 453.190 0.000 453.470 4.000 ;
=======
        RECT 272.410 0.000 272.690 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 462.390 0.000 462.670 4.000 ;
=======
        RECT 277.930 0.000 278.210 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 471.590 0.000 471.870 4.000 ;
=======
        RECT 283.450 0.000 283.730 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 480.790 0.000 481.070 4.000 ;
=======
        RECT 288.970 0.000 289.250 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 489.990 0.000 490.270 4.000 ;
=======
        RECT 294.490 0.000 294.770 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 498.730 0.000 499.010 4.000 ;
=======
        RECT 300.010 0.000 300.290 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 334.970 0.000 335.250 4.000 ;
=======
        RECT 201.110 0.000 201.390 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 507.930 0.000 508.210 4.000 ;
=======
        RECT 305.070 0.000 305.350 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 517.130 0.000 517.410 4.000 ;
=======
        RECT 310.590 0.000 310.870 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 526.330 0.000 526.610 4.000 ;
=======
        RECT 316.110 0.000 316.390 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 535.530 0.000 535.810 4.000 ;
=======
        RECT 321.630 0.000 321.910 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 544.270 0.000 544.550 4.000 ;
=======
        RECT 327.150 0.000 327.430 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 553.470 0.000 553.750 4.000 ;
=======
        RECT 332.670 0.000 332.950 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 562.670 0.000 562.950 4.000 ;
=======
        RECT 338.190 0.000 338.470 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 571.870 0.000 572.150 4.000 ;
=======
        RECT 343.710 0.000 343.990 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 580.610 0.000 580.890 4.000 ;
=======
        RECT 349.230 0.000 349.510 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 589.810 0.000 590.090 4.000 ;
=======
        RECT 354.750 0.000 355.030 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 344.170 0.000 344.450 4.000 ;
=======
        RECT 206.630 0.000 206.910 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 599.010 0.000 599.290 4.000 ;
=======
        RECT 360.270 0.000 360.550 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 608.210 0.000 608.490 4.000 ;
=======
        RECT 365.330 0.000 365.610 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 617.410 0.000 617.690 4.000 ;
=======
        RECT 370.850 0.000 371.130 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 626.150 0.000 626.430 4.000 ;
=======
        RECT 376.370 0.000 376.650 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 635.350 0.000 635.630 4.000 ;
=======
        RECT 381.890 0.000 382.170 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 644.550 0.000 644.830 4.000 ;
=======
        RECT 387.410 0.000 387.690 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 653.750 0.000 654.030 4.000 ;
=======
        RECT 392.930 0.000 393.210 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 662.950 0.000 663.230 4.000 ;
=======
        RECT 398.450 0.000 398.730 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 671.690 0.000 671.970 4.000 ;
=======
        RECT 403.970 0.000 404.250 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 680.890 0.000 681.170 4.000 ;
=======
        RECT 409.490 0.000 409.770 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 353.370 0.000 353.650 4.000 ;
=======
        RECT 212.150 0.000 212.430 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 690.090 0.000 690.370 4.000 ;
=======
        RECT 415.010 0.000 415.290 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 699.290 0.000 699.570 4.000 ;
=======
        RECT 420.530 0.000 420.810 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 708.490 0.000 708.770 4.000 ;
=======
        RECT 425.590 0.000 425.870 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 717.230 0.000 717.510 4.000 ;
=======
        RECT 431.110 0.000 431.390 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 726.430 0.000 726.710 4.000 ;
=======
        RECT 436.630 0.000 436.910 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 735.630 0.000 735.910 4.000 ;
=======
        RECT 442.150 0.000 442.430 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 744.830 0.000 745.110 4.000 ;
=======
        RECT 447.670 0.000 447.950 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 753.570 0.000 753.850 4.000 ;
=======
        RECT 453.190 0.000 453.470 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 762.770 0.000 763.050 4.000 ;
=======
        RECT 458.710 0.000 458.990 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 771.970 0.000 772.250 4.000 ;
=======
        RECT 464.230 0.000 464.510 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 362.570 0.000 362.850 4.000 ;
=======
        RECT 217.670 0.000 217.950 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 781.170 0.000 781.450 4.000 ;
=======
        RECT 469.750 0.000 470.030 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 790.370 0.000 790.650 4.000 ;
=======
        RECT 475.270 0.000 475.550 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 799.110 0.000 799.390 4.000 ;
=======
        RECT 480.330 0.000 480.610 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 808.310 0.000 808.590 4.000 ;
=======
        RECT 485.850 0.000 486.130 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 817.510 0.000 817.790 4.000 ;
=======
        RECT 491.370 0.000 491.650 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 826.710 0.000 826.990 4.000 ;
=======
        RECT 496.890 0.000 497.170 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 835.910 0.000 836.190 4.000 ;
=======
        RECT 502.410 0.000 502.690 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 844.650 0.000 844.930 4.000 ;
=======
        RECT 507.930 0.000 508.210 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 853.850 0.000 854.130 4.000 ;
=======
        RECT 513.450 0.000 513.730 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 863.050 0.000 863.330 4.000 ;
=======
        RECT 518.970 0.000 519.250 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 371.310 0.000 371.590 4.000 ;
=======
        RECT 223.190 0.000 223.470 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 872.250 0.000 872.530 4.000 ;
=======
        RECT 524.490 0.000 524.770 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 881.450 0.000 881.730 4.000 ;
=======
        RECT 530.010 0.000 530.290 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 890.190 0.000 890.470 4.000 ;
=======
        RECT 535.530 0.000 535.810 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 899.390 0.000 899.670 4.000 ;
=======
        RECT 540.590 0.000 540.870 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 908.590 0.000 908.870 4.000 ;
=======
        RECT 546.110 0.000 546.390 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 917.790 0.000 918.070 4.000 ;
=======
        RECT 551.630 0.000 551.910 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 926.990 0.000 927.270 4.000 ;
=======
        RECT 557.150 0.000 557.430 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 935.730 0.000 936.010 4.000 ;
=======
        RECT 562.670 0.000 562.950 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 944.930 0.000 945.210 4.000 ;
=======
        RECT 568.190 0.000 568.470 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 954.130 0.000 954.410 4.000 ;
=======
        RECT 573.710 0.000 573.990 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 380.510 0.000 380.790 4.000 ;
=======
        RECT 228.710 0.000 228.990 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 963.330 0.000 963.610 4.000 ;
=======
        RECT 579.230 0.000 579.510 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 972.070 0.000 972.350 4.000 ;
=======
        RECT 584.750 0.000 585.030 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 981.270 0.000 981.550 4.000 ;
=======
        RECT 590.270 0.000 590.550 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 990.470 0.000 990.750 4.000 ;
=======
        RECT 595.790 0.000 596.070 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 999.670 0.000 999.950 4.000 ;
=======
        RECT 600.850 0.000 601.130 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1008.870 0.000 1009.150 4.000 ;
=======
        RECT 606.370 0.000 606.650 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1017.610 0.000 1017.890 4.000 ;
=======
        RECT 611.890 0.000 612.170 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1026.810 0.000 1027.090 4.000 ;
=======
        RECT 617.410 0.000 617.690 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1036.010 0.000 1036.290 4.000 ;
=======
        RECT 622.930 0.000 623.210 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1045.210 0.000 1045.490 4.000 ;
=======
        RECT 628.450 0.000 628.730 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 389.710 0.000 389.990 4.000 ;
=======
        RECT 234.230 0.000 234.510 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1054.410 0.000 1054.690 4.000 ;
=======
        RECT 633.970 0.000 634.250 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1063.150 0.000 1063.430 4.000 ;
=======
        RECT 639.490 0.000 639.770 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1072.350 0.000 1072.630 4.000 ;
=======
        RECT 645.010 0.000 645.290 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1081.550 0.000 1081.830 4.000 ;
=======
        RECT 650.530 0.000 650.810 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1090.750 0.000 1091.030 4.000 ;
=======
        RECT 656.050 0.000 656.330 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1099.950 0.000 1100.230 4.000 ;
=======
        RECT 661.110 0.000 661.390 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1108.690 0.000 1108.970 4.000 ;
=======
        RECT 666.630 0.000 666.910 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1117.890 0.000 1118.170 4.000 ;
=======
        RECT 672.150 0.000 672.430 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1127.090 0.000 1127.370 4.000 ;
=======
        RECT 677.670 0.000 677.950 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1136.290 0.000 1136.570 4.000 ;
=======
        RECT 683.190 0.000 683.470 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 398.910 0.000 399.190 4.000 ;
=======
        RECT 239.750 0.000 240.030 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1145.030 0.000 1145.310 4.000 ;
=======
        RECT 688.710 0.000 688.990 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1154.230 0.000 1154.510 4.000 ;
=======
        RECT 694.230 0.000 694.510 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1163.430 0.000 1163.710 4.000 ;
=======
        RECT 699.750 0.000 700.030 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1172.630 0.000 1172.910 4.000 ;
=======
        RECT 705.270 0.000 705.550 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1181.830 0.000 1182.110 4.000 ;
=======
        RECT 710.790 0.000 711.070 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1190.570 0.000 1190.850 4.000 ;
=======
        RECT 716.310 0.000 716.590 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1199.770 0.000 1200.050 4.000 ;
=======
        RECT 721.370 0.000 721.650 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1208.970 0.000 1209.250 4.000 ;
=======
        RECT 726.890 0.000 727.170 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1218.170 0.000 1218.450 4.000 ;
=======
        RECT 732.410 0.000 732.690 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1227.370 0.000 1227.650 4.000 ;
=======
        RECT 737.930 0.000 738.210 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 407.650 0.000 407.930 4.000 ;
=======
        RECT 244.810 0.000 245.090 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 328.990 0.000 329.270 4.000 ;
=======
        RECT 197.430 0.000 197.710 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1239.330 0.000 1239.610 4.000 ;
=======
        RECT 745.290 0.000 745.570 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1248.530 0.000 1248.810 4.000 ;
=======
        RECT 750.810 0.000 751.090 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1257.730 0.000 1258.010 4.000 ;
=======
        RECT 756.330 0.000 756.610 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1266.470 0.000 1266.750 4.000 ;
=======
        RECT 761.850 0.000 762.130 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1275.670 0.000 1275.950 4.000 ;
=======
        RECT 767.370 0.000 767.650 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1284.870 0.000 1285.150 4.000 ;
=======
        RECT 772.890 0.000 773.170 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1294.070 0.000 1294.350 4.000 ;
=======
        RECT 778.410 0.000 778.690 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1303.270 0.000 1303.550 4.000 ;
=======
        RECT 783.470 0.000 783.750 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1312.010 0.000 1312.290 4.000 ;
=======
        RECT 788.990 0.000 789.270 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1321.210 0.000 1321.490 4.000 ;
=======
        RECT 794.510 0.000 794.790 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 420.070 0.000 420.350 4.000 ;
=======
        RECT 252.170 0.000 252.450 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1330.410 0.000 1330.690 4.000 ;
=======
        RECT 800.030 0.000 800.310 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1339.610 0.000 1339.890 4.000 ;
=======
        RECT 805.550 0.000 805.830 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1348.350 0.000 1348.630 4.000 ;
=======
        RECT 811.070 0.000 811.350 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1357.550 0.000 1357.830 4.000 ;
=======
        RECT 816.590 0.000 816.870 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1366.750 0.000 1367.030 4.000 ;
=======
        RECT 822.110 0.000 822.390 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1375.950 0.000 1376.230 4.000 ;
=======
        RECT 827.630 0.000 827.910 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1385.150 0.000 1385.430 4.000 ;
=======
        RECT 833.150 0.000 833.430 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1393.890 0.000 1394.170 4.000 ;
=======
        RECT 838.670 0.000 838.950 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1403.090 0.000 1403.370 4.000 ;
=======
        RECT 843.730 0.000 844.010 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1412.290 0.000 1412.570 4.000 ;
=======
        RECT 849.250 0.000 849.530 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 429.270 0.000 429.550 4.000 ;
=======
        RECT 257.690 0.000 257.970 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1421.490 0.000 1421.770 4.000 ;
=======
        RECT 854.770 0.000 855.050 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1430.690 0.000 1430.970 4.000 ;
=======
        RECT 860.290 0.000 860.570 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1439.430 0.000 1439.710 4.000 ;
=======
        RECT 865.810 0.000 866.090 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1448.630 0.000 1448.910 4.000 ;
=======
        RECT 871.330 0.000 871.610 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1457.830 0.000 1458.110 4.000 ;
=======
        RECT 876.850 0.000 877.130 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1467.030 0.000 1467.310 4.000 ;
=======
        RECT 882.370 0.000 882.650 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1476.230 0.000 1476.510 4.000 ;
=======
        RECT 887.890 0.000 888.170 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1484.970 0.000 1485.250 4.000 ;
=======
        RECT 893.410 0.000 893.690 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 438.010 0.000 438.290 4.000 ;
=======
        RECT 263.210 0.000 263.490 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 447.210 0.000 447.490 4.000 ;
=======
        RECT 268.730 0.000 269.010 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 456.410 0.000 456.690 4.000 ;
=======
        RECT 274.250 0.000 274.530 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 465.610 0.000 465.890 4.000 ;
=======
        RECT 279.770 0.000 280.050 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 474.810 0.000 475.090 4.000 ;
=======
        RECT 285.290 0.000 285.570 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 483.550 0.000 483.830 4.000 ;
=======
        RECT 290.810 0.000 291.090 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 492.750 0.000 493.030 4.000 ;
=======
        RECT 296.330 0.000 296.610 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 501.950 0.000 502.230 4.000 ;
=======
        RECT 301.390 0.000 301.670 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 338.190 0.000 338.470 4.000 ;
=======
        RECT 202.950 0.000 203.230 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 511.150 0.000 511.430 4.000 ;
=======
        RECT 306.910 0.000 307.190 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 520.350 0.000 520.630 4.000 ;
=======
        RECT 312.430 0.000 312.710 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 529.090 0.000 529.370 4.000 ;
=======
        RECT 317.950 0.000 318.230 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 538.290 0.000 538.570 4.000 ;
=======
        RECT 323.470 0.000 323.750 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 547.490 0.000 547.770 4.000 ;
=======
        RECT 328.990 0.000 329.270 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 556.690 0.000 556.970 4.000 ;
=======
        RECT 334.510 0.000 334.790 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 565.430 0.000 565.710 4.000 ;
=======
        RECT 340.030 0.000 340.310 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 574.630 0.000 574.910 4.000 ;
=======
        RECT 345.550 0.000 345.830 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 583.830 0.000 584.110 4.000 ;
=======
        RECT 351.070 0.000 351.350 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 593.030 0.000 593.310 4.000 ;
=======
        RECT 356.590 0.000 356.870 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 347.390 0.000 347.670 4.000 ;
=======
        RECT 208.470 0.000 208.750 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 602.230 0.000 602.510 4.000 ;
=======
        RECT 361.650 0.000 361.930 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 610.970 0.000 611.250 4.000 ;
=======
        RECT 367.170 0.000 367.450 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 620.170 0.000 620.450 4.000 ;
=======
        RECT 372.690 0.000 372.970 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 629.370 0.000 629.650 4.000 ;
=======
        RECT 378.210 0.000 378.490 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 638.570 0.000 638.850 4.000 ;
=======
        RECT 383.730 0.000 384.010 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 647.770 0.000 648.050 4.000 ;
=======
        RECT 389.250 0.000 389.530 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 656.510 0.000 656.790 4.000 ;
=======
        RECT 394.770 0.000 395.050 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 665.710 0.000 665.990 4.000 ;
=======
        RECT 400.290 0.000 400.570 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 674.910 0.000 675.190 4.000 ;
=======
        RECT 405.810 0.000 406.090 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 684.110 0.000 684.390 4.000 ;
=======
        RECT 411.330 0.000 411.610 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 356.130 0.000 356.410 4.000 ;
=======
        RECT 213.990 0.000 214.270 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 693.310 0.000 693.590 4.000 ;
=======
        RECT 416.850 0.000 417.130 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 702.050 0.000 702.330 4.000 ;
=======
        RECT 421.910 0.000 422.190 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 711.250 0.000 711.530 4.000 ;
=======
        RECT 427.430 0.000 427.710 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 720.450 0.000 720.730 4.000 ;
=======
        RECT 432.950 0.000 433.230 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 729.650 0.000 729.930 4.000 ;
=======
        RECT 438.470 0.000 438.750 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 738.850 0.000 739.130 4.000 ;
=======
        RECT 443.990 0.000 444.270 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 747.590 0.000 747.870 4.000 ;
=======
        RECT 449.510 0.000 449.790 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 756.790 0.000 757.070 4.000 ;
=======
        RECT 455.030 0.000 455.310 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 765.990 0.000 766.270 4.000 ;
=======
        RECT 460.550 0.000 460.830 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 775.190 0.000 775.470 4.000 ;
=======
        RECT 466.070 0.000 466.350 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 365.330 0.000 365.610 4.000 ;
=======
        RECT 219.510 0.000 219.790 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 783.930 0.000 784.210 4.000 ;
=======
        RECT 471.590 0.000 471.870 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 793.130 0.000 793.410 4.000 ;
=======
        RECT 477.110 0.000 477.390 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 802.330 0.000 802.610 4.000 ;
=======
        RECT 482.170 0.000 482.450 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 811.530 0.000 811.810 4.000 ;
=======
        RECT 487.690 0.000 487.970 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 820.730 0.000 821.010 4.000 ;
=======
        RECT 493.210 0.000 493.490 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 829.470 0.000 829.750 4.000 ;
=======
        RECT 498.730 0.000 499.010 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 838.670 0.000 838.950 4.000 ;
=======
        RECT 504.250 0.000 504.530 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 847.870 0.000 848.150 4.000 ;
=======
        RECT 509.770 0.000 510.050 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 857.070 0.000 857.350 4.000 ;
=======
        RECT 515.290 0.000 515.570 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 866.270 0.000 866.550 4.000 ;
=======
        RECT 520.810 0.000 521.090 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 374.530 0.000 374.810 4.000 ;
=======
        RECT 225.030 0.000 225.310 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 875.010 0.000 875.290 4.000 ;
=======
        RECT 526.330 0.000 526.610 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 884.210 0.000 884.490 4.000 ;
=======
        RECT 531.850 0.000 532.130 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 893.410 0.000 893.690 4.000 ;
=======
        RECT 537.370 0.000 537.650 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 902.610 0.000 902.890 4.000 ;
=======
        RECT 542.430 0.000 542.710 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 911.810 0.000 912.090 4.000 ;
=======
        RECT 547.950 0.000 548.230 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 920.550 0.000 920.830 4.000 ;
=======
        RECT 553.470 0.000 553.750 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 929.750 0.000 930.030 4.000 ;
=======
        RECT 558.990 0.000 559.270 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 938.950 0.000 939.230 4.000 ;
=======
        RECT 564.510 0.000 564.790 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 948.150 0.000 948.430 4.000 ;
=======
        RECT 570.030 0.000 570.310 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 956.890 0.000 957.170 4.000 ;
=======
        RECT 575.550 0.000 575.830 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 383.730 0.000 384.010 4.000 ;
=======
        RECT 230.550 0.000 230.830 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 966.090 0.000 966.370 4.000 ;
=======
        RECT 581.070 0.000 581.350 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 975.290 0.000 975.570 4.000 ;
=======
        RECT 586.590 0.000 586.870 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 984.490 0.000 984.770 4.000 ;
=======
        RECT 592.110 0.000 592.390 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 993.690 0.000 993.970 4.000 ;
=======
        RECT 597.630 0.000 597.910 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1002.430 0.000 1002.710 4.000 ;
=======
        RECT 602.690 0.000 602.970 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1011.630 0.000 1011.910 4.000 ;
=======
        RECT 608.210 0.000 608.490 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1020.830 0.000 1021.110 4.000 ;
=======
        RECT 613.730 0.000 614.010 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1030.030 0.000 1030.310 4.000 ;
=======
        RECT 619.250 0.000 619.530 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1039.230 0.000 1039.510 4.000 ;
=======
        RECT 624.770 0.000 625.050 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1047.970 0.000 1048.250 4.000 ;
=======
        RECT 630.290 0.000 630.570 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 392.470 0.000 392.750 4.000 ;
=======
        RECT 236.070 0.000 236.350 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1057.170 0.000 1057.450 4.000 ;
=======
        RECT 635.810 0.000 636.090 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1066.370 0.000 1066.650 4.000 ;
=======
        RECT 641.330 0.000 641.610 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1075.570 0.000 1075.850 4.000 ;
=======
        RECT 646.850 0.000 647.130 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1084.770 0.000 1085.050 4.000 ;
=======
        RECT 652.370 0.000 652.650 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1093.510 0.000 1093.790 4.000 ;
=======
        RECT 657.890 0.000 658.170 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1102.710 0.000 1102.990 4.000 ;
=======
        RECT 662.950 0.000 663.230 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1111.910 0.000 1112.190 4.000 ;
=======
        RECT 668.470 0.000 668.750 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1121.110 0.000 1121.390 4.000 ;
=======
        RECT 673.990 0.000 674.270 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1129.850 0.000 1130.130 4.000 ;
=======
        RECT 679.510 0.000 679.790 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1139.050 0.000 1139.330 4.000 ;
=======
        RECT 685.030 0.000 685.310 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 401.670 0.000 401.950 4.000 ;
=======
        RECT 241.130 0.000 241.410 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1148.250 0.000 1148.530 4.000 ;
=======
        RECT 690.550 0.000 690.830 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1157.450 0.000 1157.730 4.000 ;
=======
        RECT 696.070 0.000 696.350 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1166.650 0.000 1166.930 4.000 ;
=======
        RECT 701.590 0.000 701.870 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1175.390 0.000 1175.670 4.000 ;
=======
        RECT 707.110 0.000 707.390 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1184.590 0.000 1184.870 4.000 ;
=======
        RECT 712.630 0.000 712.910 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1193.790 0.000 1194.070 4.000 ;
=======
        RECT 718.150 0.000 718.430 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1202.990 0.000 1203.270 4.000 ;
=======
        RECT 723.210 0.000 723.490 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1212.190 0.000 1212.470 4.000 ;
=======
        RECT 728.730 0.000 729.010 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1220.930 0.000 1221.210 4.000 ;
=======
        RECT 734.250 0.000 734.530 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 1230.130 0.000 1230.410 4.000 ;
=======
        RECT 739.770 0.000 740.050 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 410.870 0.000 411.150 4.000 ;
    END
  END la_oenb[9]
  PIN user_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1488.190 0.000 1488.470 4.000 ;
    END
  END user_clk
=======
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END la_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 122.450 0.000 122.730 4.000 ;
=======
        RECT 73.230 0.000 73.510 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 131.650 0.000 131.930 4.000 ;
=======
        RECT 78.750 0.000 79.030 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 140.850 0.000 141.130 4.000 ;
=======
        RECT 84.270 0.000 84.550 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 150.050 0.000 150.330 4.000 ;
=======
        RECT 89.790 0.000 90.070 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 159.250 0.000 159.530 4.000 ;
=======
        RECT 95.310 0.000 95.590 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 167.990 0.000 168.270 4.000 ;
=======
        RECT 100.830 0.000 101.110 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 177.190 0.000 177.470 4.000 ;
=======
        RECT 106.350 0.000 106.630 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 186.390 0.000 186.670 4.000 ;
=======
        RECT 111.870 0.000 112.150 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 195.590 0.000 195.870 4.000 ;
=======
        RECT 117.390 0.000 117.670 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 204.330 0.000 204.610 4.000 ;
=======
        RECT 122.450 0.000 122.730 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 213.530 0.000 213.810 4.000 ;
=======
        RECT 127.970 0.000 128.250 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 222.730 0.000 223.010 4.000 ;
=======
        RECT 133.490 0.000 133.770 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 231.930 0.000 232.210 4.000 ;
=======
        RECT 139.010 0.000 139.290 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 241.130 0.000 241.410 4.000 ;
=======
        RECT 144.530 0.000 144.810 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 249.870 0.000 250.150 4.000 ;
=======
        RECT 150.050 0.000 150.330 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 259.070 0.000 259.350 4.000 ;
=======
        RECT 155.570 0.000 155.850 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 268.270 0.000 268.550 4.000 ;
=======
        RECT 161.090 0.000 161.370 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 277.470 0.000 277.750 4.000 ;
=======
        RECT 166.610 0.000 166.890 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 286.670 0.000 286.950 4.000 ;
=======
        RECT 172.130 0.000 172.410 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 295.410 0.000 295.690 4.000 ;
=======
        RECT 177.650 0.000 177.930 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 304.610 0.000 304.890 4.000 ;
=======
        RECT 182.710 0.000 182.990 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 313.810 0.000 314.090 4.000 ;
=======
        RECT 188.230 0.000 188.510 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 104.510 0.000 104.790 4.000 ;
=======
        RECT 62.190 0.000 62.470 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 113.710 0.000 113.990 4.000 ;
=======
        RECT 67.710 0.000 67.990 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 125.670 0.000 125.950 4.000 ;
=======
        RECT 75.070 0.000 75.350 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 134.870 0.000 135.150 4.000 ;
=======
        RECT 80.590 0.000 80.870 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 144.070 0.000 144.350 4.000 ;
=======
        RECT 86.110 0.000 86.390 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 152.810 0.000 153.090 4.000 ;
=======
        RECT 91.630 0.000 91.910 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 162.010 0.000 162.290 4.000 ;
=======
        RECT 97.150 0.000 97.430 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 171.210 0.000 171.490 4.000 ;
=======
        RECT 102.670 0.000 102.950 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 180.410 0.000 180.690 4.000 ;
=======
        RECT 108.190 0.000 108.470 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 189.150 0.000 189.430 4.000 ;
=======
        RECT 113.710 0.000 113.990 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 198.350 0.000 198.630 4.000 ;
=======
        RECT 119.230 0.000 119.510 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 207.550 0.000 207.830 4.000 ;
=======
        RECT 124.290 0.000 124.570 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 216.750 0.000 217.030 4.000 ;
=======
        RECT 129.810 0.000 130.090 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 225.950 0.000 226.230 4.000 ;
=======
        RECT 135.330 0.000 135.610 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 234.690 0.000 234.970 4.000 ;
=======
        RECT 140.850 0.000 141.130 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 243.890 0.000 244.170 4.000 ;
=======
        RECT 146.370 0.000 146.650 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 253.090 0.000 253.370 4.000 ;
=======
        RECT 151.890 0.000 152.170 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 262.290 0.000 262.570 4.000 ;
=======
        RECT 157.410 0.000 157.690 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 271.490 0.000 271.770 4.000 ;
=======
        RECT 162.930 0.000 163.210 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 280.230 0.000 280.510 4.000 ;
=======
        RECT 168.450 0.000 168.730 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 289.430 0.000 289.710 4.000 ;
=======
        RECT 173.970 0.000 174.250 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 298.630 0.000 298.910 4.000 ;
=======
        RECT 179.490 0.000 179.770 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 307.830 0.000 308.110 4.000 ;
=======
        RECT 184.550 0.000 184.830 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 317.030 0.000 317.310 4.000 ;
=======
        RECT 190.070 0.000 190.350 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 107.270 0.000 107.550 4.000 ;
=======
        RECT 64.030 0.000 64.310 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 116.470 0.000 116.750 4.000 ;
=======
        RECT 69.550 0.000 69.830 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 128.890 0.000 129.170 4.000 ;
=======
        RECT 76.910 0.000 77.190 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 137.630 0.000 137.910 4.000 ;
=======
        RECT 82.430 0.000 82.710 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 146.830 0.000 147.110 4.000 ;
=======
        RECT 87.950 0.000 88.230 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 156.030 0.000 156.310 4.000 ;
=======
        RECT 93.470 0.000 93.750 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 165.230 0.000 165.510 4.000 ;
=======
        RECT 98.990 0.000 99.270 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 174.430 0.000 174.710 4.000 ;
=======
        RECT 104.510 0.000 104.790 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 183.170 0.000 183.450 4.000 ;
=======
        RECT 110.030 0.000 110.310 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 192.370 0.000 192.650 4.000 ;
=======
        RECT 115.550 0.000 115.830 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 201.570 0.000 201.850 4.000 ;
=======
        RECT 120.610 0.000 120.890 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 210.770 0.000 211.050 4.000 ;
=======
        RECT 126.130 0.000 126.410 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 219.510 0.000 219.790 4.000 ;
=======
        RECT 131.650 0.000 131.930 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 228.710 0.000 228.990 4.000 ;
=======
        RECT 137.170 0.000 137.450 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 237.910 0.000 238.190 4.000 ;
=======
        RECT 142.690 0.000 142.970 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 247.110 0.000 247.390 4.000 ;
=======
        RECT 148.210 0.000 148.490 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 256.310 0.000 256.590 4.000 ;
=======
        RECT 153.730 0.000 154.010 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 265.050 0.000 265.330 4.000 ;
=======
        RECT 159.250 0.000 159.530 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 274.250 0.000 274.530 4.000 ;
=======
        RECT 164.770 0.000 165.050 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 283.450 0.000 283.730 4.000 ;
=======
        RECT 170.290 0.000 170.570 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 292.650 0.000 292.930 4.000 ;
=======
        RECT 175.810 0.000 176.090 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 301.850 0.000 302.130 4.000 ;
=======
        RECT 180.870 0.000 181.150 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 310.590 0.000 310.870 4.000 ;
=======
        RECT 186.390 0.000 186.670 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 319.790 0.000 320.070 4.000 ;
=======
        RECT 191.910 0.000 192.190 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 101.290 0.000 101.570 4.000 ;
=======
        RECT 60.350 0.000 60.630 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 110.490 0.000 110.770 4.000 ;
=======
        RECT 65.870 0.000 66.150 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 119.690 0.000 119.970 4.000 ;
=======
        RECT 71.390 0.000 71.670 4.000 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END wbs_we_i
<<<<<<< HEAD
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1477.200 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1477.200 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1477.200 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1477.200 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1477.200 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1477.200 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1477.200 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1477.200 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1477.200 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1477.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1477.200 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1477.200 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1477.200 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1477.200 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1477.200 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1477.200 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1477.200 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1477.200 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1477.200 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1477.200 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1406.740 10.880 1408.340 1476.960 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1253.140 10.880 1254.740 1476.960 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1099.540 10.880 1101.140 1476.960 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 945.940 10.880 947.540 1476.960 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 792.340 10.880 793.940 1476.960 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 1476.960 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 1476.960 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 1476.960 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 1476.960 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 1476.960 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1329.940 10.880 1331.540 1476.960 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1176.340 10.880 1177.940 1476.960 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1022.740 10.880 1024.340 1476.960 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 869.140 10.880 870.740 1476.960 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 715.540 10.880 717.140 1476.960 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 1476.960 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 1476.960 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 1476.960 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 1476.960 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1410.040 10.880 1411.640 1476.960 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1256.440 10.880 1258.040 1476.960 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1102.840 10.880 1104.440 1476.960 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 949.240 10.880 950.840 1476.960 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 795.640 10.880 797.240 1476.960 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 642.040 10.880 643.640 1476.960 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.440 10.880 490.040 1476.960 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 1476.960 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 1476.960 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 1476.960 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1333.240 10.880 1334.840 1476.960 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1179.640 10.880 1181.240 1476.960 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1026.040 10.880 1027.640 1476.960 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 872.440 10.880 874.040 1476.960 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 718.840 10.880 720.440 1476.960 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 565.240 10.880 566.840 1476.960 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.640 10.880 413.240 1476.960 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 1476.960 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 1476.960 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1413.340 10.880 1414.940 1476.960 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1259.740 10.880 1261.340 1476.960 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1106.140 10.880 1107.740 1476.960 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 952.540 10.880 954.140 1476.960 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 798.940 10.880 800.540 1476.960 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 645.340 10.880 646.940 1476.960 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.740 10.880 493.340 1476.960 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 1476.960 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 1476.960 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 1476.960 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1336.540 10.880 1338.140 1476.960 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1182.940 10.880 1184.540 1476.960 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1029.340 10.880 1030.940 1476.960 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 875.740 10.880 877.340 1476.960 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 722.140 10.880 723.740 1476.960 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.540 10.880 570.140 1476.960 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.940 10.880 416.540 1476.960 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 1476.960 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 1476.960 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 5.525 1484.420 1477.045 ;
      LAYER met1 ;
        RECT 1.450 4.800 1488.490 1477.200 ;
      LAYER met2 ;
        RECT 1.480 1485.720 5.790 1486.000 ;
        RECT 6.630 1485.720 18.210 1486.000 ;
        RECT 19.050 1485.720 31.090 1486.000 ;
        RECT 31.930 1485.720 43.970 1486.000 ;
        RECT 44.810 1485.720 56.850 1486.000 ;
        RECT 57.690 1485.720 69.730 1486.000 ;
        RECT 70.570 1485.720 82.610 1486.000 ;
        RECT 83.450 1485.720 95.490 1486.000 ;
        RECT 96.330 1485.720 108.370 1486.000 ;
        RECT 109.210 1485.720 121.250 1486.000 ;
        RECT 122.090 1485.720 134.130 1486.000 ;
        RECT 134.970 1485.720 147.010 1486.000 ;
        RECT 147.850 1485.720 159.890 1486.000 ;
        RECT 160.730 1485.720 172.310 1486.000 ;
        RECT 173.150 1485.720 185.190 1486.000 ;
        RECT 186.030 1485.720 198.070 1486.000 ;
        RECT 198.910 1485.720 210.950 1486.000 ;
        RECT 211.790 1485.720 223.830 1486.000 ;
        RECT 224.670 1485.720 236.710 1486.000 ;
        RECT 237.550 1485.720 249.590 1486.000 ;
        RECT 250.430 1485.720 262.470 1486.000 ;
        RECT 263.310 1485.720 275.350 1486.000 ;
        RECT 276.190 1485.720 288.230 1486.000 ;
        RECT 289.070 1485.720 301.110 1486.000 ;
        RECT 301.950 1485.720 313.990 1486.000 ;
        RECT 314.830 1485.720 326.870 1486.000 ;
        RECT 327.710 1485.720 339.290 1486.000 ;
        RECT 340.130 1485.720 352.170 1486.000 ;
        RECT 353.010 1485.720 365.050 1486.000 ;
        RECT 365.890 1485.720 377.930 1486.000 ;
        RECT 378.770 1485.720 390.810 1486.000 ;
        RECT 391.650 1485.720 403.690 1486.000 ;
        RECT 404.530 1485.720 416.570 1486.000 ;
        RECT 417.410 1485.720 429.450 1486.000 ;
        RECT 430.290 1485.720 442.330 1486.000 ;
        RECT 443.170 1485.720 455.210 1486.000 ;
        RECT 456.050 1485.720 468.090 1486.000 ;
        RECT 468.930 1485.720 480.970 1486.000 ;
        RECT 481.810 1485.720 493.850 1486.000 ;
        RECT 494.690 1485.720 506.270 1486.000 ;
        RECT 507.110 1485.720 519.150 1486.000 ;
        RECT 519.990 1485.720 532.030 1486.000 ;
        RECT 532.870 1485.720 544.910 1486.000 ;
        RECT 545.750 1485.720 557.790 1486.000 ;
        RECT 558.630 1485.720 570.670 1486.000 ;
        RECT 571.510 1485.720 583.550 1486.000 ;
        RECT 584.390 1485.720 596.430 1486.000 ;
        RECT 597.270 1485.720 609.310 1486.000 ;
        RECT 610.150 1485.720 622.190 1486.000 ;
        RECT 623.030 1485.720 635.070 1486.000 ;
        RECT 635.910 1485.720 647.950 1486.000 ;
        RECT 648.790 1485.720 660.830 1486.000 ;
        RECT 661.670 1485.720 673.250 1486.000 ;
        RECT 674.090 1485.720 686.130 1486.000 ;
        RECT 686.970 1485.720 699.010 1486.000 ;
        RECT 699.850 1485.720 711.890 1486.000 ;
        RECT 712.730 1485.720 724.770 1486.000 ;
        RECT 725.610 1485.720 737.650 1486.000 ;
        RECT 738.490 1485.720 750.530 1486.000 ;
        RECT 751.370 1485.720 763.410 1486.000 ;
        RECT 764.250 1485.720 776.290 1486.000 ;
        RECT 777.130 1485.720 789.170 1486.000 ;
        RECT 790.010 1485.720 802.050 1486.000 ;
        RECT 802.890 1485.720 814.930 1486.000 ;
        RECT 815.770 1485.720 827.810 1486.000 ;
        RECT 828.650 1485.720 840.230 1486.000 ;
        RECT 841.070 1485.720 853.110 1486.000 ;
        RECT 853.950 1485.720 865.990 1486.000 ;
        RECT 866.830 1485.720 878.870 1486.000 ;
        RECT 879.710 1485.720 891.750 1486.000 ;
        RECT 892.590 1485.720 904.630 1486.000 ;
        RECT 905.470 1485.720 917.510 1486.000 ;
        RECT 918.350 1485.720 930.390 1486.000 ;
        RECT 931.230 1485.720 943.270 1486.000 ;
        RECT 944.110 1485.720 956.150 1486.000 ;
        RECT 956.990 1485.720 969.030 1486.000 ;
        RECT 969.870 1485.720 981.910 1486.000 ;
        RECT 982.750 1485.720 994.790 1486.000 ;
        RECT 995.630 1485.720 1007.210 1486.000 ;
        RECT 1008.050 1485.720 1020.090 1486.000 ;
        RECT 1020.930 1485.720 1032.970 1486.000 ;
        RECT 1033.810 1485.720 1045.850 1486.000 ;
        RECT 1046.690 1485.720 1058.730 1486.000 ;
        RECT 1059.570 1485.720 1071.610 1486.000 ;
        RECT 1072.450 1485.720 1084.490 1486.000 ;
        RECT 1085.330 1485.720 1097.370 1486.000 ;
        RECT 1098.210 1485.720 1110.250 1486.000 ;
        RECT 1111.090 1485.720 1123.130 1486.000 ;
        RECT 1123.970 1485.720 1136.010 1486.000 ;
        RECT 1136.850 1485.720 1148.890 1486.000 ;
        RECT 1149.730 1485.720 1161.770 1486.000 ;
        RECT 1162.610 1485.720 1174.190 1486.000 ;
        RECT 1175.030 1485.720 1187.070 1486.000 ;
        RECT 1187.910 1485.720 1199.950 1486.000 ;
        RECT 1200.790 1485.720 1212.830 1486.000 ;
        RECT 1213.670 1485.720 1225.710 1486.000 ;
        RECT 1226.550 1485.720 1238.590 1486.000 ;
        RECT 1239.430 1485.720 1251.470 1486.000 ;
        RECT 1252.310 1485.720 1264.350 1486.000 ;
        RECT 1265.190 1485.720 1277.230 1486.000 ;
        RECT 1278.070 1485.720 1290.110 1486.000 ;
        RECT 1290.950 1485.720 1302.990 1486.000 ;
        RECT 1303.830 1485.720 1315.870 1486.000 ;
        RECT 1316.710 1485.720 1328.750 1486.000 ;
        RECT 1329.590 1485.720 1341.170 1486.000 ;
        RECT 1342.010 1485.720 1354.050 1486.000 ;
        RECT 1354.890 1485.720 1366.930 1486.000 ;
        RECT 1367.770 1485.720 1379.810 1486.000 ;
        RECT 1380.650 1485.720 1392.690 1486.000 ;
        RECT 1393.530 1485.720 1405.570 1486.000 ;
        RECT 1406.410 1485.720 1418.450 1486.000 ;
        RECT 1419.290 1485.720 1431.330 1486.000 ;
        RECT 1432.170 1485.720 1444.210 1486.000 ;
        RECT 1445.050 1485.720 1457.090 1486.000 ;
        RECT 1457.930 1485.720 1469.970 1486.000 ;
        RECT 1470.810 1485.720 1482.850 1486.000 ;
        RECT 1483.690 1485.720 1488.460 1486.000 ;
        RECT 1.480 4.280 1488.460 1485.720 ;
        RECT 2.030 4.000 3.950 4.280 ;
        RECT 4.790 4.000 7.170 4.280 ;
        RECT 8.010 4.000 9.930 4.280 ;
        RECT 10.770 4.000 13.150 4.280 ;
        RECT 13.990 4.000 15.910 4.280 ;
        RECT 16.750 4.000 19.130 4.280 ;
        RECT 19.970 4.000 22.350 4.280 ;
        RECT 23.190 4.000 25.110 4.280 ;
        RECT 25.950 4.000 28.330 4.280 ;
        RECT 29.170 4.000 31.090 4.280 ;
        RECT 31.930 4.000 34.310 4.280 ;
        RECT 35.150 4.000 37.530 4.280 ;
        RECT 38.370 4.000 40.290 4.280 ;
        RECT 41.130 4.000 43.510 4.280 ;
        RECT 44.350 4.000 46.270 4.280 ;
        RECT 47.110 4.000 49.490 4.280 ;
        RECT 50.330 4.000 52.710 4.280 ;
        RECT 53.550 4.000 55.470 4.280 ;
        RECT 56.310 4.000 58.690 4.280 ;
        RECT 59.530 4.000 61.450 4.280 ;
        RECT 62.290 4.000 64.670 4.280 ;
        RECT 65.510 4.000 67.890 4.280 ;
        RECT 68.730 4.000 70.650 4.280 ;
        RECT 71.490 4.000 73.870 4.280 ;
        RECT 74.710 4.000 76.630 4.280 ;
        RECT 77.470 4.000 79.850 4.280 ;
        RECT 80.690 4.000 83.070 4.280 ;
        RECT 83.910 4.000 85.830 4.280 ;
        RECT 86.670 4.000 89.050 4.280 ;
        RECT 89.890 4.000 91.810 4.280 ;
        RECT 92.650 4.000 95.030 4.280 ;
        RECT 95.870 4.000 98.250 4.280 ;
        RECT 99.090 4.000 101.010 4.280 ;
        RECT 101.850 4.000 104.230 4.280 ;
        RECT 105.070 4.000 106.990 4.280 ;
        RECT 107.830 4.000 110.210 4.280 ;
        RECT 111.050 4.000 113.430 4.280 ;
        RECT 114.270 4.000 116.190 4.280 ;
        RECT 117.030 4.000 119.410 4.280 ;
        RECT 120.250 4.000 122.170 4.280 ;
        RECT 123.010 4.000 125.390 4.280 ;
        RECT 126.230 4.000 128.610 4.280 ;
        RECT 129.450 4.000 131.370 4.280 ;
        RECT 132.210 4.000 134.590 4.280 ;
        RECT 135.430 4.000 137.350 4.280 ;
        RECT 138.190 4.000 140.570 4.280 ;
        RECT 141.410 4.000 143.790 4.280 ;
        RECT 144.630 4.000 146.550 4.280 ;
        RECT 147.390 4.000 149.770 4.280 ;
        RECT 150.610 4.000 152.530 4.280 ;
        RECT 153.370 4.000 155.750 4.280 ;
        RECT 156.590 4.000 158.970 4.280 ;
        RECT 159.810 4.000 161.730 4.280 ;
        RECT 162.570 4.000 164.950 4.280 ;
        RECT 165.790 4.000 167.710 4.280 ;
        RECT 168.550 4.000 170.930 4.280 ;
        RECT 171.770 4.000 174.150 4.280 ;
        RECT 174.990 4.000 176.910 4.280 ;
        RECT 177.750 4.000 180.130 4.280 ;
        RECT 180.970 4.000 182.890 4.280 ;
        RECT 183.730 4.000 186.110 4.280 ;
        RECT 186.950 4.000 188.870 4.280 ;
        RECT 189.710 4.000 192.090 4.280 ;
        RECT 192.930 4.000 195.310 4.280 ;
        RECT 196.150 4.000 198.070 4.280 ;
        RECT 198.910 4.000 201.290 4.280 ;
        RECT 202.130 4.000 204.050 4.280 ;
        RECT 204.890 4.000 207.270 4.280 ;
        RECT 208.110 4.000 210.490 4.280 ;
        RECT 211.330 4.000 213.250 4.280 ;
        RECT 214.090 4.000 216.470 4.280 ;
        RECT 217.310 4.000 219.230 4.280 ;
        RECT 220.070 4.000 222.450 4.280 ;
        RECT 223.290 4.000 225.670 4.280 ;
        RECT 226.510 4.000 228.430 4.280 ;
        RECT 229.270 4.000 231.650 4.280 ;
        RECT 232.490 4.000 234.410 4.280 ;
        RECT 235.250 4.000 237.630 4.280 ;
        RECT 238.470 4.000 240.850 4.280 ;
        RECT 241.690 4.000 243.610 4.280 ;
        RECT 244.450 4.000 246.830 4.280 ;
        RECT 247.670 4.000 249.590 4.280 ;
        RECT 250.430 4.000 252.810 4.280 ;
        RECT 253.650 4.000 256.030 4.280 ;
        RECT 256.870 4.000 258.790 4.280 ;
        RECT 259.630 4.000 262.010 4.280 ;
        RECT 262.850 4.000 264.770 4.280 ;
        RECT 265.610 4.000 267.990 4.280 ;
        RECT 268.830 4.000 271.210 4.280 ;
        RECT 272.050 4.000 273.970 4.280 ;
        RECT 274.810 4.000 277.190 4.280 ;
        RECT 278.030 4.000 279.950 4.280 ;
        RECT 280.790 4.000 283.170 4.280 ;
        RECT 284.010 4.000 286.390 4.280 ;
        RECT 287.230 4.000 289.150 4.280 ;
        RECT 289.990 4.000 292.370 4.280 ;
        RECT 293.210 4.000 295.130 4.280 ;
        RECT 295.970 4.000 298.350 4.280 ;
        RECT 299.190 4.000 301.570 4.280 ;
        RECT 302.410 4.000 304.330 4.280 ;
        RECT 305.170 4.000 307.550 4.280 ;
        RECT 308.390 4.000 310.310 4.280 ;
        RECT 311.150 4.000 313.530 4.280 ;
        RECT 314.370 4.000 316.750 4.280 ;
        RECT 317.590 4.000 319.510 4.280 ;
        RECT 320.350 4.000 322.730 4.280 ;
        RECT 323.570 4.000 325.490 4.280 ;
        RECT 326.330 4.000 328.710 4.280 ;
        RECT 329.550 4.000 331.930 4.280 ;
        RECT 332.770 4.000 334.690 4.280 ;
        RECT 335.530 4.000 337.910 4.280 ;
        RECT 338.750 4.000 340.670 4.280 ;
        RECT 341.510 4.000 343.890 4.280 ;
        RECT 344.730 4.000 347.110 4.280 ;
        RECT 347.950 4.000 349.870 4.280 ;
        RECT 350.710 4.000 353.090 4.280 ;
        RECT 353.930 4.000 355.850 4.280 ;
        RECT 356.690 4.000 359.070 4.280 ;
        RECT 359.910 4.000 362.290 4.280 ;
        RECT 363.130 4.000 365.050 4.280 ;
        RECT 365.890 4.000 368.270 4.280 ;
        RECT 369.110 4.000 371.030 4.280 ;
        RECT 371.870 4.000 374.250 4.280 ;
        RECT 375.090 4.000 377.010 4.280 ;
        RECT 377.850 4.000 380.230 4.280 ;
        RECT 381.070 4.000 383.450 4.280 ;
        RECT 384.290 4.000 386.210 4.280 ;
        RECT 387.050 4.000 389.430 4.280 ;
        RECT 390.270 4.000 392.190 4.280 ;
        RECT 393.030 4.000 395.410 4.280 ;
        RECT 396.250 4.000 398.630 4.280 ;
        RECT 399.470 4.000 401.390 4.280 ;
        RECT 402.230 4.000 404.610 4.280 ;
        RECT 405.450 4.000 407.370 4.280 ;
        RECT 408.210 4.000 410.590 4.280 ;
        RECT 411.430 4.000 413.810 4.280 ;
        RECT 414.650 4.000 416.570 4.280 ;
        RECT 417.410 4.000 419.790 4.280 ;
        RECT 420.630 4.000 422.550 4.280 ;
        RECT 423.390 4.000 425.770 4.280 ;
        RECT 426.610 4.000 428.990 4.280 ;
        RECT 429.830 4.000 431.750 4.280 ;
        RECT 432.590 4.000 434.970 4.280 ;
        RECT 435.810 4.000 437.730 4.280 ;
        RECT 438.570 4.000 440.950 4.280 ;
        RECT 441.790 4.000 444.170 4.280 ;
        RECT 445.010 4.000 446.930 4.280 ;
        RECT 447.770 4.000 450.150 4.280 ;
        RECT 450.990 4.000 452.910 4.280 ;
        RECT 453.750 4.000 456.130 4.280 ;
        RECT 456.970 4.000 459.350 4.280 ;
        RECT 460.190 4.000 462.110 4.280 ;
        RECT 462.950 4.000 465.330 4.280 ;
        RECT 466.170 4.000 468.090 4.280 ;
        RECT 468.930 4.000 471.310 4.280 ;
        RECT 472.150 4.000 474.530 4.280 ;
        RECT 475.370 4.000 477.290 4.280 ;
        RECT 478.130 4.000 480.510 4.280 ;
        RECT 481.350 4.000 483.270 4.280 ;
        RECT 484.110 4.000 486.490 4.280 ;
        RECT 487.330 4.000 489.710 4.280 ;
        RECT 490.550 4.000 492.470 4.280 ;
        RECT 493.310 4.000 495.690 4.280 ;
        RECT 496.530 4.000 498.450 4.280 ;
        RECT 499.290 4.000 501.670 4.280 ;
        RECT 502.510 4.000 504.890 4.280 ;
        RECT 505.730 4.000 507.650 4.280 ;
        RECT 508.490 4.000 510.870 4.280 ;
        RECT 511.710 4.000 513.630 4.280 ;
        RECT 514.470 4.000 516.850 4.280 ;
        RECT 517.690 4.000 520.070 4.280 ;
        RECT 520.910 4.000 522.830 4.280 ;
        RECT 523.670 4.000 526.050 4.280 ;
        RECT 526.890 4.000 528.810 4.280 ;
        RECT 529.650 4.000 532.030 4.280 ;
        RECT 532.870 4.000 535.250 4.280 ;
        RECT 536.090 4.000 538.010 4.280 ;
        RECT 538.850 4.000 541.230 4.280 ;
        RECT 542.070 4.000 543.990 4.280 ;
        RECT 544.830 4.000 547.210 4.280 ;
        RECT 548.050 4.000 550.430 4.280 ;
        RECT 551.270 4.000 553.190 4.280 ;
        RECT 554.030 4.000 556.410 4.280 ;
        RECT 557.250 4.000 559.170 4.280 ;
        RECT 560.010 4.000 562.390 4.280 ;
        RECT 563.230 4.000 565.150 4.280 ;
        RECT 565.990 4.000 568.370 4.280 ;
        RECT 569.210 4.000 571.590 4.280 ;
        RECT 572.430 4.000 574.350 4.280 ;
        RECT 575.190 4.000 577.570 4.280 ;
        RECT 578.410 4.000 580.330 4.280 ;
        RECT 581.170 4.000 583.550 4.280 ;
        RECT 584.390 4.000 586.770 4.280 ;
        RECT 587.610 4.000 589.530 4.280 ;
        RECT 590.370 4.000 592.750 4.280 ;
        RECT 593.590 4.000 595.510 4.280 ;
        RECT 596.350 4.000 598.730 4.280 ;
        RECT 599.570 4.000 601.950 4.280 ;
        RECT 602.790 4.000 604.710 4.280 ;
        RECT 605.550 4.000 607.930 4.280 ;
        RECT 608.770 4.000 610.690 4.280 ;
        RECT 611.530 4.000 613.910 4.280 ;
        RECT 614.750 4.000 617.130 4.280 ;
        RECT 617.970 4.000 619.890 4.280 ;
        RECT 620.730 4.000 623.110 4.280 ;
        RECT 623.950 4.000 625.870 4.280 ;
        RECT 626.710 4.000 629.090 4.280 ;
        RECT 629.930 4.000 632.310 4.280 ;
        RECT 633.150 4.000 635.070 4.280 ;
        RECT 635.910 4.000 638.290 4.280 ;
        RECT 639.130 4.000 641.050 4.280 ;
        RECT 641.890 4.000 644.270 4.280 ;
        RECT 645.110 4.000 647.490 4.280 ;
        RECT 648.330 4.000 650.250 4.280 ;
        RECT 651.090 4.000 653.470 4.280 ;
        RECT 654.310 4.000 656.230 4.280 ;
        RECT 657.070 4.000 659.450 4.280 ;
        RECT 660.290 4.000 662.670 4.280 ;
        RECT 663.510 4.000 665.430 4.280 ;
        RECT 666.270 4.000 668.650 4.280 ;
        RECT 669.490 4.000 671.410 4.280 ;
        RECT 672.250 4.000 674.630 4.280 ;
        RECT 675.470 4.000 677.850 4.280 ;
        RECT 678.690 4.000 680.610 4.280 ;
        RECT 681.450 4.000 683.830 4.280 ;
        RECT 684.670 4.000 686.590 4.280 ;
        RECT 687.430 4.000 689.810 4.280 ;
        RECT 690.650 4.000 693.030 4.280 ;
        RECT 693.870 4.000 695.790 4.280 ;
        RECT 696.630 4.000 699.010 4.280 ;
        RECT 699.850 4.000 701.770 4.280 ;
        RECT 702.610 4.000 704.990 4.280 ;
        RECT 705.830 4.000 708.210 4.280 ;
        RECT 709.050 4.000 710.970 4.280 ;
        RECT 711.810 4.000 714.190 4.280 ;
        RECT 715.030 4.000 716.950 4.280 ;
        RECT 717.790 4.000 720.170 4.280 ;
        RECT 721.010 4.000 723.390 4.280 ;
        RECT 724.230 4.000 726.150 4.280 ;
        RECT 726.990 4.000 729.370 4.280 ;
        RECT 730.210 4.000 732.130 4.280 ;
        RECT 732.970 4.000 735.350 4.280 ;
        RECT 736.190 4.000 738.570 4.280 ;
        RECT 739.410 4.000 741.330 4.280 ;
        RECT 742.170 4.000 744.550 4.280 ;
        RECT 745.390 4.000 747.310 4.280 ;
        RECT 748.150 4.000 750.530 4.280 ;
        RECT 751.370 4.000 753.290 4.280 ;
        RECT 754.130 4.000 756.510 4.280 ;
        RECT 757.350 4.000 759.730 4.280 ;
        RECT 760.570 4.000 762.490 4.280 ;
        RECT 763.330 4.000 765.710 4.280 ;
        RECT 766.550 4.000 768.470 4.280 ;
        RECT 769.310 4.000 771.690 4.280 ;
        RECT 772.530 4.000 774.910 4.280 ;
        RECT 775.750 4.000 777.670 4.280 ;
        RECT 778.510 4.000 780.890 4.280 ;
        RECT 781.730 4.000 783.650 4.280 ;
        RECT 784.490 4.000 786.870 4.280 ;
        RECT 787.710 4.000 790.090 4.280 ;
        RECT 790.930 4.000 792.850 4.280 ;
        RECT 793.690 4.000 796.070 4.280 ;
        RECT 796.910 4.000 798.830 4.280 ;
        RECT 799.670 4.000 802.050 4.280 ;
        RECT 802.890 4.000 805.270 4.280 ;
        RECT 806.110 4.000 808.030 4.280 ;
        RECT 808.870 4.000 811.250 4.280 ;
        RECT 812.090 4.000 814.010 4.280 ;
        RECT 814.850 4.000 817.230 4.280 ;
        RECT 818.070 4.000 820.450 4.280 ;
        RECT 821.290 4.000 823.210 4.280 ;
        RECT 824.050 4.000 826.430 4.280 ;
        RECT 827.270 4.000 829.190 4.280 ;
        RECT 830.030 4.000 832.410 4.280 ;
        RECT 833.250 4.000 835.630 4.280 ;
        RECT 836.470 4.000 838.390 4.280 ;
        RECT 839.230 4.000 841.610 4.280 ;
        RECT 842.450 4.000 844.370 4.280 ;
        RECT 845.210 4.000 847.590 4.280 ;
        RECT 848.430 4.000 850.810 4.280 ;
        RECT 851.650 4.000 853.570 4.280 ;
        RECT 854.410 4.000 856.790 4.280 ;
        RECT 857.630 4.000 859.550 4.280 ;
        RECT 860.390 4.000 862.770 4.280 ;
        RECT 863.610 4.000 865.990 4.280 ;
        RECT 866.830 4.000 868.750 4.280 ;
        RECT 869.590 4.000 871.970 4.280 ;
        RECT 872.810 4.000 874.730 4.280 ;
        RECT 875.570 4.000 877.950 4.280 ;
        RECT 878.790 4.000 881.170 4.280 ;
        RECT 882.010 4.000 883.930 4.280 ;
        RECT 884.770 4.000 887.150 4.280 ;
        RECT 887.990 4.000 889.910 4.280 ;
        RECT 890.750 4.000 893.130 4.280 ;
        RECT 893.970 4.000 896.350 4.280 ;
        RECT 897.190 4.000 899.110 4.280 ;
        RECT 899.950 4.000 902.330 4.280 ;
        RECT 903.170 4.000 905.090 4.280 ;
        RECT 905.930 4.000 908.310 4.280 ;
        RECT 909.150 4.000 911.530 4.280 ;
        RECT 912.370 4.000 914.290 4.280 ;
        RECT 915.130 4.000 917.510 4.280 ;
        RECT 918.350 4.000 920.270 4.280 ;
        RECT 921.110 4.000 923.490 4.280 ;
        RECT 924.330 4.000 926.710 4.280 ;
        RECT 927.550 4.000 929.470 4.280 ;
        RECT 930.310 4.000 932.690 4.280 ;
        RECT 933.530 4.000 935.450 4.280 ;
        RECT 936.290 4.000 938.670 4.280 ;
        RECT 939.510 4.000 941.430 4.280 ;
        RECT 942.270 4.000 944.650 4.280 ;
        RECT 945.490 4.000 947.870 4.280 ;
        RECT 948.710 4.000 950.630 4.280 ;
        RECT 951.470 4.000 953.850 4.280 ;
        RECT 954.690 4.000 956.610 4.280 ;
        RECT 957.450 4.000 959.830 4.280 ;
        RECT 960.670 4.000 963.050 4.280 ;
        RECT 963.890 4.000 965.810 4.280 ;
        RECT 966.650 4.000 969.030 4.280 ;
        RECT 969.870 4.000 971.790 4.280 ;
        RECT 972.630 4.000 975.010 4.280 ;
        RECT 975.850 4.000 978.230 4.280 ;
        RECT 979.070 4.000 980.990 4.280 ;
        RECT 981.830 4.000 984.210 4.280 ;
        RECT 985.050 4.000 986.970 4.280 ;
        RECT 987.810 4.000 990.190 4.280 ;
        RECT 991.030 4.000 993.410 4.280 ;
        RECT 994.250 4.000 996.170 4.280 ;
        RECT 997.010 4.000 999.390 4.280 ;
        RECT 1000.230 4.000 1002.150 4.280 ;
        RECT 1002.990 4.000 1005.370 4.280 ;
        RECT 1006.210 4.000 1008.590 4.280 ;
        RECT 1009.430 4.000 1011.350 4.280 ;
        RECT 1012.190 4.000 1014.570 4.280 ;
        RECT 1015.410 4.000 1017.330 4.280 ;
        RECT 1018.170 4.000 1020.550 4.280 ;
        RECT 1021.390 4.000 1023.770 4.280 ;
        RECT 1024.610 4.000 1026.530 4.280 ;
        RECT 1027.370 4.000 1029.750 4.280 ;
        RECT 1030.590 4.000 1032.510 4.280 ;
        RECT 1033.350 4.000 1035.730 4.280 ;
        RECT 1036.570 4.000 1038.950 4.280 ;
        RECT 1039.790 4.000 1041.710 4.280 ;
        RECT 1042.550 4.000 1044.930 4.280 ;
        RECT 1045.770 4.000 1047.690 4.280 ;
        RECT 1048.530 4.000 1050.910 4.280 ;
        RECT 1051.750 4.000 1054.130 4.280 ;
        RECT 1054.970 4.000 1056.890 4.280 ;
        RECT 1057.730 4.000 1060.110 4.280 ;
        RECT 1060.950 4.000 1062.870 4.280 ;
        RECT 1063.710 4.000 1066.090 4.280 ;
        RECT 1066.930 4.000 1069.310 4.280 ;
        RECT 1070.150 4.000 1072.070 4.280 ;
        RECT 1072.910 4.000 1075.290 4.280 ;
        RECT 1076.130 4.000 1078.050 4.280 ;
        RECT 1078.890 4.000 1081.270 4.280 ;
        RECT 1082.110 4.000 1084.490 4.280 ;
        RECT 1085.330 4.000 1087.250 4.280 ;
        RECT 1088.090 4.000 1090.470 4.280 ;
        RECT 1091.310 4.000 1093.230 4.280 ;
        RECT 1094.070 4.000 1096.450 4.280 ;
        RECT 1097.290 4.000 1099.670 4.280 ;
        RECT 1100.510 4.000 1102.430 4.280 ;
        RECT 1103.270 4.000 1105.650 4.280 ;
        RECT 1106.490 4.000 1108.410 4.280 ;
        RECT 1109.250 4.000 1111.630 4.280 ;
        RECT 1112.470 4.000 1114.850 4.280 ;
        RECT 1115.690 4.000 1117.610 4.280 ;
        RECT 1118.450 4.000 1120.830 4.280 ;
        RECT 1121.670 4.000 1123.590 4.280 ;
        RECT 1124.430 4.000 1126.810 4.280 ;
        RECT 1127.650 4.000 1129.570 4.280 ;
        RECT 1130.410 4.000 1132.790 4.280 ;
        RECT 1133.630 4.000 1136.010 4.280 ;
        RECT 1136.850 4.000 1138.770 4.280 ;
        RECT 1139.610 4.000 1141.990 4.280 ;
        RECT 1142.830 4.000 1144.750 4.280 ;
        RECT 1145.590 4.000 1147.970 4.280 ;
        RECT 1148.810 4.000 1151.190 4.280 ;
        RECT 1152.030 4.000 1153.950 4.280 ;
        RECT 1154.790 4.000 1157.170 4.280 ;
        RECT 1158.010 4.000 1159.930 4.280 ;
        RECT 1160.770 4.000 1163.150 4.280 ;
        RECT 1163.990 4.000 1166.370 4.280 ;
        RECT 1167.210 4.000 1169.130 4.280 ;
        RECT 1169.970 4.000 1172.350 4.280 ;
        RECT 1173.190 4.000 1175.110 4.280 ;
        RECT 1175.950 4.000 1178.330 4.280 ;
        RECT 1179.170 4.000 1181.550 4.280 ;
        RECT 1182.390 4.000 1184.310 4.280 ;
        RECT 1185.150 4.000 1187.530 4.280 ;
        RECT 1188.370 4.000 1190.290 4.280 ;
        RECT 1191.130 4.000 1193.510 4.280 ;
        RECT 1194.350 4.000 1196.730 4.280 ;
        RECT 1197.570 4.000 1199.490 4.280 ;
        RECT 1200.330 4.000 1202.710 4.280 ;
        RECT 1203.550 4.000 1205.470 4.280 ;
        RECT 1206.310 4.000 1208.690 4.280 ;
        RECT 1209.530 4.000 1211.910 4.280 ;
        RECT 1212.750 4.000 1214.670 4.280 ;
        RECT 1215.510 4.000 1217.890 4.280 ;
        RECT 1218.730 4.000 1220.650 4.280 ;
        RECT 1221.490 4.000 1223.870 4.280 ;
        RECT 1224.710 4.000 1227.090 4.280 ;
        RECT 1227.930 4.000 1229.850 4.280 ;
        RECT 1230.690 4.000 1233.070 4.280 ;
        RECT 1233.910 4.000 1235.830 4.280 ;
        RECT 1236.670 4.000 1239.050 4.280 ;
        RECT 1239.890 4.000 1242.270 4.280 ;
        RECT 1243.110 4.000 1245.030 4.280 ;
        RECT 1245.870 4.000 1248.250 4.280 ;
        RECT 1249.090 4.000 1251.010 4.280 ;
        RECT 1251.850 4.000 1254.230 4.280 ;
        RECT 1255.070 4.000 1257.450 4.280 ;
        RECT 1258.290 4.000 1260.210 4.280 ;
        RECT 1261.050 4.000 1263.430 4.280 ;
        RECT 1264.270 4.000 1266.190 4.280 ;
        RECT 1267.030 4.000 1269.410 4.280 ;
        RECT 1270.250 4.000 1272.630 4.280 ;
        RECT 1273.470 4.000 1275.390 4.280 ;
        RECT 1276.230 4.000 1278.610 4.280 ;
        RECT 1279.450 4.000 1281.370 4.280 ;
        RECT 1282.210 4.000 1284.590 4.280 ;
        RECT 1285.430 4.000 1287.810 4.280 ;
        RECT 1288.650 4.000 1290.570 4.280 ;
        RECT 1291.410 4.000 1293.790 4.280 ;
        RECT 1294.630 4.000 1296.550 4.280 ;
        RECT 1297.390 4.000 1299.770 4.280 ;
        RECT 1300.610 4.000 1302.990 4.280 ;
        RECT 1303.830 4.000 1305.750 4.280 ;
        RECT 1306.590 4.000 1308.970 4.280 ;
        RECT 1309.810 4.000 1311.730 4.280 ;
        RECT 1312.570 4.000 1314.950 4.280 ;
        RECT 1315.790 4.000 1317.710 4.280 ;
        RECT 1318.550 4.000 1320.930 4.280 ;
        RECT 1321.770 4.000 1324.150 4.280 ;
        RECT 1324.990 4.000 1326.910 4.280 ;
        RECT 1327.750 4.000 1330.130 4.280 ;
        RECT 1330.970 4.000 1332.890 4.280 ;
        RECT 1333.730 4.000 1336.110 4.280 ;
        RECT 1336.950 4.000 1339.330 4.280 ;
        RECT 1340.170 4.000 1342.090 4.280 ;
        RECT 1342.930 4.000 1345.310 4.280 ;
        RECT 1346.150 4.000 1348.070 4.280 ;
        RECT 1348.910 4.000 1351.290 4.280 ;
        RECT 1352.130 4.000 1354.510 4.280 ;
        RECT 1355.350 4.000 1357.270 4.280 ;
        RECT 1358.110 4.000 1360.490 4.280 ;
        RECT 1361.330 4.000 1363.250 4.280 ;
        RECT 1364.090 4.000 1366.470 4.280 ;
        RECT 1367.310 4.000 1369.690 4.280 ;
        RECT 1370.530 4.000 1372.450 4.280 ;
        RECT 1373.290 4.000 1375.670 4.280 ;
        RECT 1376.510 4.000 1378.430 4.280 ;
        RECT 1379.270 4.000 1381.650 4.280 ;
        RECT 1382.490 4.000 1384.870 4.280 ;
        RECT 1385.710 4.000 1387.630 4.280 ;
        RECT 1388.470 4.000 1390.850 4.280 ;
        RECT 1391.690 4.000 1393.610 4.280 ;
        RECT 1394.450 4.000 1396.830 4.280 ;
        RECT 1397.670 4.000 1400.050 4.280 ;
        RECT 1400.890 4.000 1402.810 4.280 ;
        RECT 1403.650 4.000 1406.030 4.280 ;
        RECT 1406.870 4.000 1408.790 4.280 ;
        RECT 1409.630 4.000 1412.010 4.280 ;
        RECT 1412.850 4.000 1415.230 4.280 ;
        RECT 1416.070 4.000 1417.990 4.280 ;
        RECT 1418.830 4.000 1421.210 4.280 ;
        RECT 1422.050 4.000 1423.970 4.280 ;
        RECT 1424.810 4.000 1427.190 4.280 ;
        RECT 1428.030 4.000 1430.410 4.280 ;
        RECT 1431.250 4.000 1433.170 4.280 ;
        RECT 1434.010 4.000 1436.390 4.280 ;
        RECT 1437.230 4.000 1439.150 4.280 ;
        RECT 1439.990 4.000 1442.370 4.280 ;
        RECT 1443.210 4.000 1445.590 4.280 ;
        RECT 1446.430 4.000 1448.350 4.280 ;
        RECT 1449.190 4.000 1451.570 4.280 ;
        RECT 1452.410 4.000 1454.330 4.280 ;
        RECT 1455.170 4.000 1457.550 4.280 ;
        RECT 1458.390 4.000 1460.770 4.280 ;
        RECT 1461.610 4.000 1463.530 4.280 ;
        RECT 1464.370 4.000 1466.750 4.280 ;
        RECT 1467.590 4.000 1469.510 4.280 ;
        RECT 1470.350 4.000 1472.730 4.280 ;
        RECT 1473.570 4.000 1475.950 4.280 ;
        RECT 1476.790 4.000 1478.710 4.280 ;
        RECT 1479.550 4.000 1481.930 4.280 ;
        RECT 1482.770 4.000 1484.690 4.280 ;
        RECT 1485.530 4.000 1487.910 4.280 ;
      LAYER met3 ;
        RECT 4.000 745.640 1483.435 1477.125 ;
        RECT 4.400 744.240 1483.435 745.640 ;
        RECT 4.000 6.975 1483.435 744.240 ;
      LAYER met4 ;
        RECT 23.295 15.815 23.940 1448.225 ;
        RECT 26.340 15.815 27.240 1448.225 ;
        RECT 29.640 15.815 30.540 1448.225 ;
        RECT 32.940 15.815 97.440 1448.225 ;
        RECT 99.840 15.815 100.740 1448.225 ;
        RECT 103.140 15.815 104.040 1448.225 ;
        RECT 106.440 15.815 107.340 1448.225 ;
        RECT 109.740 15.815 174.240 1448.225 ;
        RECT 176.640 15.815 177.540 1448.225 ;
        RECT 179.940 15.815 180.840 1448.225 ;
        RECT 183.240 15.815 184.140 1448.225 ;
        RECT 186.540 15.815 251.040 1448.225 ;
        RECT 253.440 15.815 254.340 1448.225 ;
        RECT 256.740 15.815 257.640 1448.225 ;
        RECT 260.040 15.815 260.940 1448.225 ;
        RECT 263.340 15.815 327.840 1448.225 ;
        RECT 330.240 15.815 331.140 1448.225 ;
        RECT 333.540 15.815 334.440 1448.225 ;
        RECT 336.840 15.815 337.740 1448.225 ;
        RECT 340.140 15.815 404.640 1448.225 ;
        RECT 407.040 15.815 407.940 1448.225 ;
        RECT 410.340 15.815 411.240 1448.225 ;
        RECT 413.640 15.815 414.540 1448.225 ;
        RECT 416.940 15.815 481.440 1448.225 ;
        RECT 483.840 15.815 484.740 1448.225 ;
        RECT 487.140 15.815 488.040 1448.225 ;
        RECT 490.440 15.815 491.340 1448.225 ;
        RECT 493.740 15.815 558.240 1448.225 ;
        RECT 560.640 15.815 561.540 1448.225 ;
        RECT 563.940 15.815 564.840 1448.225 ;
        RECT 567.240 15.815 568.140 1448.225 ;
        RECT 570.540 15.815 635.040 1448.225 ;
        RECT 637.440 15.815 638.340 1448.225 ;
        RECT 640.740 15.815 641.640 1448.225 ;
        RECT 644.040 15.815 644.940 1448.225 ;
        RECT 647.340 15.815 711.840 1448.225 ;
        RECT 714.240 15.815 715.140 1448.225 ;
        RECT 717.540 15.815 718.440 1448.225 ;
        RECT 720.840 15.815 721.740 1448.225 ;
        RECT 724.140 15.815 788.640 1448.225 ;
        RECT 791.040 15.815 791.940 1448.225 ;
        RECT 794.340 15.815 795.240 1448.225 ;
        RECT 797.640 15.815 798.540 1448.225 ;
        RECT 800.940 15.815 865.440 1448.225 ;
        RECT 867.840 15.815 868.740 1448.225 ;
        RECT 871.140 15.815 872.040 1448.225 ;
        RECT 874.440 15.815 875.340 1448.225 ;
        RECT 877.740 15.815 942.240 1448.225 ;
        RECT 944.640 15.815 945.540 1448.225 ;
        RECT 947.940 15.815 948.840 1448.225 ;
        RECT 951.240 15.815 952.140 1448.225 ;
        RECT 954.540 15.815 1019.040 1448.225 ;
        RECT 1021.440 15.815 1022.340 1448.225 ;
        RECT 1024.740 15.815 1025.640 1448.225 ;
        RECT 1028.040 15.815 1028.940 1448.225 ;
        RECT 1031.340 15.815 1095.840 1448.225 ;
        RECT 1098.240 15.815 1099.140 1448.225 ;
        RECT 1101.540 15.815 1102.440 1448.225 ;
        RECT 1104.840 15.815 1105.740 1448.225 ;
        RECT 1108.140 15.815 1172.640 1448.225 ;
        RECT 1175.040 15.815 1175.940 1448.225 ;
        RECT 1178.340 15.815 1179.240 1448.225 ;
        RECT 1181.640 15.815 1182.540 1448.225 ;
        RECT 1184.940 15.815 1249.440 1448.225 ;
        RECT 1251.840 15.815 1252.740 1448.225 ;
        RECT 1255.140 15.815 1256.040 1448.225 ;
        RECT 1258.440 15.815 1259.340 1448.225 ;
        RECT 1261.740 15.815 1326.240 1448.225 ;
        RECT 1328.640 15.815 1329.540 1448.225 ;
        RECT 1331.940 15.815 1332.840 1448.225 ;
        RECT 1335.240 15.815 1336.140 1448.225 ;
        RECT 1338.540 15.815 1403.040 1448.225 ;
        RECT 1405.440 15.815 1406.340 1448.225 ;
        RECT 1408.740 15.815 1409.640 1448.225 ;
        RECT 1412.040 15.815 1412.940 1448.225 ;
        RECT 1415.340 15.815 1441.345 1448.225 ;
=======
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 1.910 0.040 899.230 587.760 ;
      LAYER met2 ;
        RECT 0.090 595.720 3.490 596.770 ;
        RECT 4.330 595.720 11.310 596.770 ;
        RECT 12.150 595.720 19.130 596.770 ;
        RECT 19.970 595.720 26.950 596.770 ;
        RECT 27.790 595.720 34.770 596.770 ;
        RECT 35.610 595.720 42.590 596.770 ;
        RECT 43.430 595.720 50.870 596.770 ;
        RECT 51.710 595.720 58.690 596.770 ;
        RECT 59.530 595.720 66.510 596.770 ;
        RECT 67.350 595.720 74.330 596.770 ;
        RECT 75.170 595.720 82.150 596.770 ;
        RECT 82.990 595.720 89.970 596.770 ;
        RECT 90.810 595.720 98.250 596.770 ;
        RECT 99.090 595.720 106.070 596.770 ;
        RECT 106.910 595.720 113.890 596.770 ;
        RECT 114.730 595.720 121.710 596.770 ;
        RECT 122.550 595.720 129.530 596.770 ;
        RECT 130.370 595.720 137.350 596.770 ;
        RECT 138.190 595.720 145.630 596.770 ;
        RECT 146.470 595.720 153.450 596.770 ;
        RECT 154.290 595.720 161.270 596.770 ;
        RECT 162.110 595.720 169.090 596.770 ;
        RECT 169.930 595.720 176.910 596.770 ;
        RECT 177.750 595.720 184.730 596.770 ;
        RECT 185.570 595.720 193.010 596.770 ;
        RECT 193.850 595.720 200.830 596.770 ;
        RECT 201.670 595.720 208.650 596.770 ;
        RECT 209.490 595.720 216.470 596.770 ;
        RECT 217.310 595.720 224.290 596.770 ;
        RECT 225.130 595.720 232.110 596.770 ;
        RECT 232.950 595.720 240.390 596.770 ;
        RECT 241.230 595.720 248.210 596.770 ;
        RECT 249.050 595.720 256.030 596.770 ;
        RECT 256.870 595.720 263.850 596.770 ;
        RECT 264.690 595.720 271.670 596.770 ;
        RECT 272.510 595.720 279.490 596.770 ;
        RECT 280.330 595.720 287.770 596.770 ;
        RECT 288.610 595.720 295.590 596.770 ;
        RECT 296.430 595.720 303.410 596.770 ;
        RECT 304.250 595.720 311.230 596.770 ;
        RECT 312.070 595.720 319.050 596.770 ;
        RECT 319.890 595.720 326.870 596.770 ;
        RECT 327.710 595.720 335.150 596.770 ;
        RECT 335.990 595.720 342.970 596.770 ;
        RECT 343.810 595.720 350.790 596.770 ;
        RECT 351.630 595.720 358.610 596.770 ;
        RECT 359.450 595.720 366.430 596.770 ;
        RECT 367.270 595.720 374.250 596.770 ;
        RECT 375.090 595.720 382.530 596.770 ;
        RECT 383.370 595.720 390.350 596.770 ;
        RECT 391.190 595.720 398.170 596.770 ;
        RECT 399.010 595.720 405.990 596.770 ;
        RECT 406.830 595.720 413.810 596.770 ;
        RECT 414.650 595.720 421.630 596.770 ;
        RECT 422.470 595.720 429.910 596.770 ;
        RECT 430.750 595.720 437.730 596.770 ;
        RECT 438.570 595.720 445.550 596.770 ;
        RECT 446.390 595.720 453.370 596.770 ;
        RECT 454.210 595.720 461.190 596.770 ;
        RECT 462.030 595.720 469.010 596.770 ;
        RECT 469.850 595.720 477.290 596.770 ;
        RECT 478.130 595.720 485.110 596.770 ;
        RECT 485.950 595.720 492.930 596.770 ;
        RECT 493.770 595.720 500.750 596.770 ;
        RECT 501.590 595.720 508.570 596.770 ;
        RECT 509.410 595.720 516.390 596.770 ;
        RECT 517.230 595.720 524.670 596.770 ;
        RECT 525.510 595.720 532.490 596.770 ;
        RECT 533.330 595.720 540.310 596.770 ;
        RECT 541.150 595.720 548.130 596.770 ;
        RECT 548.970 595.720 555.950 596.770 ;
        RECT 556.790 595.720 563.770 596.770 ;
        RECT 564.610 595.720 572.050 596.770 ;
        RECT 572.890 595.720 579.870 596.770 ;
        RECT 580.710 595.720 587.690 596.770 ;
        RECT 588.530 595.720 595.510 596.770 ;
        RECT 596.350 595.720 603.330 596.770 ;
        RECT 604.170 595.720 611.150 596.770 ;
        RECT 611.990 595.720 619.430 596.770 ;
        RECT 620.270 595.720 627.250 596.770 ;
        RECT 628.090 595.720 635.070 596.770 ;
        RECT 635.910 595.720 642.890 596.770 ;
        RECT 643.730 595.720 650.710 596.770 ;
        RECT 651.550 595.720 658.530 596.770 ;
        RECT 659.370 595.720 666.810 596.770 ;
        RECT 667.650 595.720 674.630 596.770 ;
        RECT 675.470 595.720 682.450 596.770 ;
        RECT 683.290 595.720 690.270 596.770 ;
        RECT 691.110 595.720 698.090 596.770 ;
        RECT 698.930 595.720 705.910 596.770 ;
        RECT 706.750 595.720 714.190 596.770 ;
        RECT 715.030 595.720 722.010 596.770 ;
        RECT 722.850 595.720 729.830 596.770 ;
        RECT 730.670 595.720 737.650 596.770 ;
        RECT 738.490 595.720 745.470 596.770 ;
        RECT 746.310 595.720 753.290 596.770 ;
        RECT 754.130 595.720 761.570 596.770 ;
        RECT 762.410 595.720 769.390 596.770 ;
        RECT 770.230 595.720 777.210 596.770 ;
        RECT 778.050 595.720 785.030 596.770 ;
        RECT 785.870 595.720 792.850 596.770 ;
        RECT 793.690 595.720 800.670 596.770 ;
        RECT 801.510 595.720 808.950 596.770 ;
        RECT 809.790 595.720 816.770 596.770 ;
        RECT 817.610 595.720 824.590 596.770 ;
        RECT 825.430 595.720 832.410 596.770 ;
        RECT 833.250 595.720 840.230 596.770 ;
        RECT 841.070 595.720 848.050 596.770 ;
        RECT 848.890 595.720 856.330 596.770 ;
        RECT 857.170 595.720 864.150 596.770 ;
        RECT 864.990 595.720 871.970 596.770 ;
        RECT 872.810 595.720 879.790 596.770 ;
        RECT 880.630 595.720 887.610 596.770 ;
        RECT 888.450 595.720 895.430 596.770 ;
        RECT 896.270 595.720 899.200 596.770 ;
        RECT 0.090 4.280 899.200 595.720 ;
        RECT 0.090 0.010 0.270 4.280 ;
        RECT 1.110 0.010 1.650 4.280 ;
        RECT 2.490 0.010 3.490 4.280 ;
        RECT 4.330 0.010 5.330 4.280 ;
        RECT 6.170 0.010 7.170 4.280 ;
        RECT 8.010 0.010 9.010 4.280 ;
        RECT 9.850 0.010 10.850 4.280 ;
        RECT 11.690 0.010 12.690 4.280 ;
        RECT 13.530 0.010 14.530 4.280 ;
        RECT 15.370 0.010 16.370 4.280 ;
        RECT 17.210 0.010 18.210 4.280 ;
        RECT 19.050 0.010 20.050 4.280 ;
        RECT 20.890 0.010 21.890 4.280 ;
        RECT 22.730 0.010 23.730 4.280 ;
        RECT 24.570 0.010 25.570 4.280 ;
        RECT 26.410 0.010 27.410 4.280 ;
        RECT 28.250 0.010 29.250 4.280 ;
        RECT 30.090 0.010 31.090 4.280 ;
        RECT 31.930 0.010 32.930 4.280 ;
        RECT 33.770 0.010 34.770 4.280 ;
        RECT 35.610 0.010 36.610 4.280 ;
        RECT 37.450 0.010 38.450 4.280 ;
        RECT 39.290 0.010 40.290 4.280 ;
        RECT 41.130 0.010 42.130 4.280 ;
        RECT 42.970 0.010 43.970 4.280 ;
        RECT 44.810 0.010 45.810 4.280 ;
        RECT 46.650 0.010 47.650 4.280 ;
        RECT 48.490 0.010 49.490 4.280 ;
        RECT 50.330 0.010 51.330 4.280 ;
        RECT 52.170 0.010 53.170 4.280 ;
        RECT 54.010 0.010 55.010 4.280 ;
        RECT 55.850 0.010 56.850 4.280 ;
        RECT 57.690 0.010 58.690 4.280 ;
        RECT 59.530 0.010 60.070 4.280 ;
        RECT 60.910 0.010 61.910 4.280 ;
        RECT 62.750 0.010 63.750 4.280 ;
        RECT 64.590 0.010 65.590 4.280 ;
        RECT 66.430 0.010 67.430 4.280 ;
        RECT 68.270 0.010 69.270 4.280 ;
        RECT 70.110 0.010 71.110 4.280 ;
        RECT 71.950 0.010 72.950 4.280 ;
        RECT 73.790 0.010 74.790 4.280 ;
        RECT 75.630 0.010 76.630 4.280 ;
        RECT 77.470 0.010 78.470 4.280 ;
        RECT 79.310 0.010 80.310 4.280 ;
        RECT 81.150 0.010 82.150 4.280 ;
        RECT 82.990 0.010 83.990 4.280 ;
        RECT 84.830 0.010 85.830 4.280 ;
        RECT 86.670 0.010 87.670 4.280 ;
        RECT 88.510 0.010 89.510 4.280 ;
        RECT 90.350 0.010 91.350 4.280 ;
        RECT 92.190 0.010 93.190 4.280 ;
        RECT 94.030 0.010 95.030 4.280 ;
        RECT 95.870 0.010 96.870 4.280 ;
        RECT 97.710 0.010 98.710 4.280 ;
        RECT 99.550 0.010 100.550 4.280 ;
        RECT 101.390 0.010 102.390 4.280 ;
        RECT 103.230 0.010 104.230 4.280 ;
        RECT 105.070 0.010 106.070 4.280 ;
        RECT 106.910 0.010 107.910 4.280 ;
        RECT 108.750 0.010 109.750 4.280 ;
        RECT 110.590 0.010 111.590 4.280 ;
        RECT 112.430 0.010 113.430 4.280 ;
        RECT 114.270 0.010 115.270 4.280 ;
        RECT 116.110 0.010 117.110 4.280 ;
        RECT 117.950 0.010 118.950 4.280 ;
        RECT 119.790 0.010 120.330 4.280 ;
        RECT 121.170 0.010 122.170 4.280 ;
        RECT 123.010 0.010 124.010 4.280 ;
        RECT 124.850 0.010 125.850 4.280 ;
        RECT 126.690 0.010 127.690 4.280 ;
        RECT 128.530 0.010 129.530 4.280 ;
        RECT 130.370 0.010 131.370 4.280 ;
        RECT 132.210 0.010 133.210 4.280 ;
        RECT 134.050 0.010 135.050 4.280 ;
        RECT 135.890 0.010 136.890 4.280 ;
        RECT 137.730 0.010 138.730 4.280 ;
        RECT 139.570 0.010 140.570 4.280 ;
        RECT 141.410 0.010 142.410 4.280 ;
        RECT 143.250 0.010 144.250 4.280 ;
        RECT 145.090 0.010 146.090 4.280 ;
        RECT 146.930 0.010 147.930 4.280 ;
        RECT 148.770 0.010 149.770 4.280 ;
        RECT 150.610 0.010 151.610 4.280 ;
        RECT 152.450 0.010 153.450 4.280 ;
        RECT 154.290 0.010 155.290 4.280 ;
        RECT 156.130 0.010 157.130 4.280 ;
        RECT 157.970 0.010 158.970 4.280 ;
        RECT 159.810 0.010 160.810 4.280 ;
        RECT 161.650 0.010 162.650 4.280 ;
        RECT 163.490 0.010 164.490 4.280 ;
        RECT 165.330 0.010 166.330 4.280 ;
        RECT 167.170 0.010 168.170 4.280 ;
        RECT 169.010 0.010 170.010 4.280 ;
        RECT 170.850 0.010 171.850 4.280 ;
        RECT 172.690 0.010 173.690 4.280 ;
        RECT 174.530 0.010 175.530 4.280 ;
        RECT 176.370 0.010 177.370 4.280 ;
        RECT 178.210 0.010 179.210 4.280 ;
        RECT 180.050 0.010 180.590 4.280 ;
        RECT 181.430 0.010 182.430 4.280 ;
        RECT 183.270 0.010 184.270 4.280 ;
        RECT 185.110 0.010 186.110 4.280 ;
        RECT 186.950 0.010 187.950 4.280 ;
        RECT 188.790 0.010 189.790 4.280 ;
        RECT 190.630 0.010 191.630 4.280 ;
        RECT 192.470 0.010 193.470 4.280 ;
        RECT 194.310 0.010 195.310 4.280 ;
        RECT 196.150 0.010 197.150 4.280 ;
        RECT 197.990 0.010 198.990 4.280 ;
        RECT 199.830 0.010 200.830 4.280 ;
        RECT 201.670 0.010 202.670 4.280 ;
        RECT 203.510 0.010 204.510 4.280 ;
        RECT 205.350 0.010 206.350 4.280 ;
        RECT 207.190 0.010 208.190 4.280 ;
        RECT 209.030 0.010 210.030 4.280 ;
        RECT 210.870 0.010 211.870 4.280 ;
        RECT 212.710 0.010 213.710 4.280 ;
        RECT 214.550 0.010 215.550 4.280 ;
        RECT 216.390 0.010 217.390 4.280 ;
        RECT 218.230 0.010 219.230 4.280 ;
        RECT 220.070 0.010 221.070 4.280 ;
        RECT 221.910 0.010 222.910 4.280 ;
        RECT 223.750 0.010 224.750 4.280 ;
        RECT 225.590 0.010 226.590 4.280 ;
        RECT 227.430 0.010 228.430 4.280 ;
        RECT 229.270 0.010 230.270 4.280 ;
        RECT 231.110 0.010 232.110 4.280 ;
        RECT 232.950 0.010 233.950 4.280 ;
        RECT 234.790 0.010 235.790 4.280 ;
        RECT 236.630 0.010 237.630 4.280 ;
        RECT 238.470 0.010 239.470 4.280 ;
        RECT 240.310 0.010 240.850 4.280 ;
        RECT 241.690 0.010 242.690 4.280 ;
        RECT 243.530 0.010 244.530 4.280 ;
        RECT 245.370 0.010 246.370 4.280 ;
        RECT 247.210 0.010 248.210 4.280 ;
        RECT 249.050 0.010 250.050 4.280 ;
        RECT 250.890 0.010 251.890 4.280 ;
        RECT 252.730 0.010 253.730 4.280 ;
        RECT 254.570 0.010 255.570 4.280 ;
        RECT 256.410 0.010 257.410 4.280 ;
        RECT 258.250 0.010 259.250 4.280 ;
        RECT 260.090 0.010 261.090 4.280 ;
        RECT 261.930 0.010 262.930 4.280 ;
        RECT 263.770 0.010 264.770 4.280 ;
        RECT 265.610 0.010 266.610 4.280 ;
        RECT 267.450 0.010 268.450 4.280 ;
        RECT 269.290 0.010 270.290 4.280 ;
        RECT 271.130 0.010 272.130 4.280 ;
        RECT 272.970 0.010 273.970 4.280 ;
        RECT 274.810 0.010 275.810 4.280 ;
        RECT 276.650 0.010 277.650 4.280 ;
        RECT 278.490 0.010 279.490 4.280 ;
        RECT 280.330 0.010 281.330 4.280 ;
        RECT 282.170 0.010 283.170 4.280 ;
        RECT 284.010 0.010 285.010 4.280 ;
        RECT 285.850 0.010 286.850 4.280 ;
        RECT 287.690 0.010 288.690 4.280 ;
        RECT 289.530 0.010 290.530 4.280 ;
        RECT 291.370 0.010 292.370 4.280 ;
        RECT 293.210 0.010 294.210 4.280 ;
        RECT 295.050 0.010 296.050 4.280 ;
        RECT 296.890 0.010 297.890 4.280 ;
        RECT 298.730 0.010 299.730 4.280 ;
        RECT 300.570 0.010 301.110 4.280 ;
        RECT 301.950 0.010 302.950 4.280 ;
        RECT 303.790 0.010 304.790 4.280 ;
        RECT 305.630 0.010 306.630 4.280 ;
        RECT 307.470 0.010 308.470 4.280 ;
        RECT 309.310 0.010 310.310 4.280 ;
        RECT 311.150 0.010 312.150 4.280 ;
        RECT 312.990 0.010 313.990 4.280 ;
        RECT 314.830 0.010 315.830 4.280 ;
        RECT 316.670 0.010 317.670 4.280 ;
        RECT 318.510 0.010 319.510 4.280 ;
        RECT 320.350 0.010 321.350 4.280 ;
        RECT 322.190 0.010 323.190 4.280 ;
        RECT 324.030 0.010 325.030 4.280 ;
        RECT 325.870 0.010 326.870 4.280 ;
        RECT 327.710 0.010 328.710 4.280 ;
        RECT 329.550 0.010 330.550 4.280 ;
        RECT 331.390 0.010 332.390 4.280 ;
        RECT 333.230 0.010 334.230 4.280 ;
        RECT 335.070 0.010 336.070 4.280 ;
        RECT 336.910 0.010 337.910 4.280 ;
        RECT 338.750 0.010 339.750 4.280 ;
        RECT 340.590 0.010 341.590 4.280 ;
        RECT 342.430 0.010 343.430 4.280 ;
        RECT 344.270 0.010 345.270 4.280 ;
        RECT 346.110 0.010 347.110 4.280 ;
        RECT 347.950 0.010 348.950 4.280 ;
        RECT 349.790 0.010 350.790 4.280 ;
        RECT 351.630 0.010 352.630 4.280 ;
        RECT 353.470 0.010 354.470 4.280 ;
        RECT 355.310 0.010 356.310 4.280 ;
        RECT 357.150 0.010 358.150 4.280 ;
        RECT 358.990 0.010 359.990 4.280 ;
        RECT 360.830 0.010 361.370 4.280 ;
        RECT 362.210 0.010 363.210 4.280 ;
        RECT 364.050 0.010 365.050 4.280 ;
        RECT 365.890 0.010 366.890 4.280 ;
        RECT 367.730 0.010 368.730 4.280 ;
        RECT 369.570 0.010 370.570 4.280 ;
        RECT 371.410 0.010 372.410 4.280 ;
        RECT 373.250 0.010 374.250 4.280 ;
        RECT 375.090 0.010 376.090 4.280 ;
        RECT 376.930 0.010 377.930 4.280 ;
        RECT 378.770 0.010 379.770 4.280 ;
        RECT 380.610 0.010 381.610 4.280 ;
        RECT 382.450 0.010 383.450 4.280 ;
        RECT 384.290 0.010 385.290 4.280 ;
        RECT 386.130 0.010 387.130 4.280 ;
        RECT 387.970 0.010 388.970 4.280 ;
        RECT 389.810 0.010 390.810 4.280 ;
        RECT 391.650 0.010 392.650 4.280 ;
        RECT 393.490 0.010 394.490 4.280 ;
        RECT 395.330 0.010 396.330 4.280 ;
        RECT 397.170 0.010 398.170 4.280 ;
        RECT 399.010 0.010 400.010 4.280 ;
        RECT 400.850 0.010 401.850 4.280 ;
        RECT 402.690 0.010 403.690 4.280 ;
        RECT 404.530 0.010 405.530 4.280 ;
        RECT 406.370 0.010 407.370 4.280 ;
        RECT 408.210 0.010 409.210 4.280 ;
        RECT 410.050 0.010 411.050 4.280 ;
        RECT 411.890 0.010 412.890 4.280 ;
        RECT 413.730 0.010 414.730 4.280 ;
        RECT 415.570 0.010 416.570 4.280 ;
        RECT 417.410 0.010 418.410 4.280 ;
        RECT 419.250 0.010 420.250 4.280 ;
        RECT 421.090 0.010 421.630 4.280 ;
        RECT 422.470 0.010 423.470 4.280 ;
        RECT 424.310 0.010 425.310 4.280 ;
        RECT 426.150 0.010 427.150 4.280 ;
        RECT 427.990 0.010 428.990 4.280 ;
        RECT 429.830 0.010 430.830 4.280 ;
        RECT 431.670 0.010 432.670 4.280 ;
        RECT 433.510 0.010 434.510 4.280 ;
        RECT 435.350 0.010 436.350 4.280 ;
        RECT 437.190 0.010 438.190 4.280 ;
        RECT 439.030 0.010 440.030 4.280 ;
        RECT 440.870 0.010 441.870 4.280 ;
        RECT 442.710 0.010 443.710 4.280 ;
        RECT 444.550 0.010 445.550 4.280 ;
        RECT 446.390 0.010 447.390 4.280 ;
        RECT 448.230 0.010 449.230 4.280 ;
        RECT 450.070 0.010 451.070 4.280 ;
        RECT 451.910 0.010 452.910 4.280 ;
        RECT 453.750 0.010 454.750 4.280 ;
        RECT 455.590 0.010 456.590 4.280 ;
        RECT 457.430 0.010 458.430 4.280 ;
        RECT 459.270 0.010 460.270 4.280 ;
        RECT 461.110 0.010 462.110 4.280 ;
        RECT 462.950 0.010 463.950 4.280 ;
        RECT 464.790 0.010 465.790 4.280 ;
        RECT 466.630 0.010 467.630 4.280 ;
        RECT 468.470 0.010 469.470 4.280 ;
        RECT 470.310 0.010 471.310 4.280 ;
        RECT 472.150 0.010 473.150 4.280 ;
        RECT 473.990 0.010 474.990 4.280 ;
        RECT 475.830 0.010 476.830 4.280 ;
        RECT 477.670 0.010 478.670 4.280 ;
        RECT 479.510 0.010 480.050 4.280 ;
        RECT 480.890 0.010 481.890 4.280 ;
        RECT 482.730 0.010 483.730 4.280 ;
        RECT 484.570 0.010 485.570 4.280 ;
        RECT 486.410 0.010 487.410 4.280 ;
        RECT 488.250 0.010 489.250 4.280 ;
        RECT 490.090 0.010 491.090 4.280 ;
        RECT 491.930 0.010 492.930 4.280 ;
        RECT 493.770 0.010 494.770 4.280 ;
        RECT 495.610 0.010 496.610 4.280 ;
        RECT 497.450 0.010 498.450 4.280 ;
        RECT 499.290 0.010 500.290 4.280 ;
        RECT 501.130 0.010 502.130 4.280 ;
        RECT 502.970 0.010 503.970 4.280 ;
        RECT 504.810 0.010 505.810 4.280 ;
        RECT 506.650 0.010 507.650 4.280 ;
        RECT 508.490 0.010 509.490 4.280 ;
        RECT 510.330 0.010 511.330 4.280 ;
        RECT 512.170 0.010 513.170 4.280 ;
        RECT 514.010 0.010 515.010 4.280 ;
        RECT 515.850 0.010 516.850 4.280 ;
        RECT 517.690 0.010 518.690 4.280 ;
        RECT 519.530 0.010 520.530 4.280 ;
        RECT 521.370 0.010 522.370 4.280 ;
        RECT 523.210 0.010 524.210 4.280 ;
        RECT 525.050 0.010 526.050 4.280 ;
        RECT 526.890 0.010 527.890 4.280 ;
        RECT 528.730 0.010 529.730 4.280 ;
        RECT 530.570 0.010 531.570 4.280 ;
        RECT 532.410 0.010 533.410 4.280 ;
        RECT 534.250 0.010 535.250 4.280 ;
        RECT 536.090 0.010 537.090 4.280 ;
        RECT 537.930 0.010 538.930 4.280 ;
        RECT 539.770 0.010 540.310 4.280 ;
        RECT 541.150 0.010 542.150 4.280 ;
        RECT 542.990 0.010 543.990 4.280 ;
        RECT 544.830 0.010 545.830 4.280 ;
        RECT 546.670 0.010 547.670 4.280 ;
        RECT 548.510 0.010 549.510 4.280 ;
        RECT 550.350 0.010 551.350 4.280 ;
        RECT 552.190 0.010 553.190 4.280 ;
        RECT 554.030 0.010 555.030 4.280 ;
        RECT 555.870 0.010 556.870 4.280 ;
        RECT 557.710 0.010 558.710 4.280 ;
        RECT 559.550 0.010 560.550 4.280 ;
        RECT 561.390 0.010 562.390 4.280 ;
        RECT 563.230 0.010 564.230 4.280 ;
        RECT 565.070 0.010 566.070 4.280 ;
        RECT 566.910 0.010 567.910 4.280 ;
        RECT 568.750 0.010 569.750 4.280 ;
        RECT 570.590 0.010 571.590 4.280 ;
        RECT 572.430 0.010 573.430 4.280 ;
        RECT 574.270 0.010 575.270 4.280 ;
        RECT 576.110 0.010 577.110 4.280 ;
        RECT 577.950 0.010 578.950 4.280 ;
        RECT 579.790 0.010 580.790 4.280 ;
        RECT 581.630 0.010 582.630 4.280 ;
        RECT 583.470 0.010 584.470 4.280 ;
        RECT 585.310 0.010 586.310 4.280 ;
        RECT 587.150 0.010 588.150 4.280 ;
        RECT 588.990 0.010 589.990 4.280 ;
        RECT 590.830 0.010 591.830 4.280 ;
        RECT 592.670 0.010 593.670 4.280 ;
        RECT 594.510 0.010 595.510 4.280 ;
        RECT 596.350 0.010 597.350 4.280 ;
        RECT 598.190 0.010 599.190 4.280 ;
        RECT 600.030 0.010 600.570 4.280 ;
        RECT 601.410 0.010 602.410 4.280 ;
        RECT 603.250 0.010 604.250 4.280 ;
        RECT 605.090 0.010 606.090 4.280 ;
        RECT 606.930 0.010 607.930 4.280 ;
        RECT 608.770 0.010 609.770 4.280 ;
        RECT 610.610 0.010 611.610 4.280 ;
        RECT 612.450 0.010 613.450 4.280 ;
        RECT 614.290 0.010 615.290 4.280 ;
        RECT 616.130 0.010 617.130 4.280 ;
        RECT 617.970 0.010 618.970 4.280 ;
        RECT 619.810 0.010 620.810 4.280 ;
        RECT 621.650 0.010 622.650 4.280 ;
        RECT 623.490 0.010 624.490 4.280 ;
        RECT 625.330 0.010 626.330 4.280 ;
        RECT 627.170 0.010 628.170 4.280 ;
        RECT 629.010 0.010 630.010 4.280 ;
        RECT 630.850 0.010 631.850 4.280 ;
        RECT 632.690 0.010 633.690 4.280 ;
        RECT 634.530 0.010 635.530 4.280 ;
        RECT 636.370 0.010 637.370 4.280 ;
        RECT 638.210 0.010 639.210 4.280 ;
        RECT 640.050 0.010 641.050 4.280 ;
        RECT 641.890 0.010 642.890 4.280 ;
        RECT 643.730 0.010 644.730 4.280 ;
        RECT 645.570 0.010 646.570 4.280 ;
        RECT 647.410 0.010 648.410 4.280 ;
        RECT 649.250 0.010 650.250 4.280 ;
        RECT 651.090 0.010 652.090 4.280 ;
        RECT 652.930 0.010 653.930 4.280 ;
        RECT 654.770 0.010 655.770 4.280 ;
        RECT 656.610 0.010 657.610 4.280 ;
        RECT 658.450 0.010 659.450 4.280 ;
        RECT 660.290 0.010 660.830 4.280 ;
        RECT 661.670 0.010 662.670 4.280 ;
        RECT 663.510 0.010 664.510 4.280 ;
        RECT 665.350 0.010 666.350 4.280 ;
        RECT 667.190 0.010 668.190 4.280 ;
        RECT 669.030 0.010 670.030 4.280 ;
        RECT 670.870 0.010 671.870 4.280 ;
        RECT 672.710 0.010 673.710 4.280 ;
        RECT 674.550 0.010 675.550 4.280 ;
        RECT 676.390 0.010 677.390 4.280 ;
        RECT 678.230 0.010 679.230 4.280 ;
        RECT 680.070 0.010 681.070 4.280 ;
        RECT 681.910 0.010 682.910 4.280 ;
        RECT 683.750 0.010 684.750 4.280 ;
        RECT 685.590 0.010 686.590 4.280 ;
        RECT 687.430 0.010 688.430 4.280 ;
        RECT 689.270 0.010 690.270 4.280 ;
        RECT 691.110 0.010 692.110 4.280 ;
        RECT 692.950 0.010 693.950 4.280 ;
        RECT 694.790 0.010 695.790 4.280 ;
        RECT 696.630 0.010 697.630 4.280 ;
        RECT 698.470 0.010 699.470 4.280 ;
        RECT 700.310 0.010 701.310 4.280 ;
        RECT 702.150 0.010 703.150 4.280 ;
        RECT 703.990 0.010 704.990 4.280 ;
        RECT 705.830 0.010 706.830 4.280 ;
        RECT 707.670 0.010 708.670 4.280 ;
        RECT 709.510 0.010 710.510 4.280 ;
        RECT 711.350 0.010 712.350 4.280 ;
        RECT 713.190 0.010 714.190 4.280 ;
        RECT 715.030 0.010 716.030 4.280 ;
        RECT 716.870 0.010 717.870 4.280 ;
        RECT 718.710 0.010 719.710 4.280 ;
        RECT 720.550 0.010 721.090 4.280 ;
        RECT 721.930 0.010 722.930 4.280 ;
        RECT 723.770 0.010 724.770 4.280 ;
        RECT 725.610 0.010 726.610 4.280 ;
        RECT 727.450 0.010 728.450 4.280 ;
        RECT 729.290 0.010 730.290 4.280 ;
        RECT 731.130 0.010 732.130 4.280 ;
        RECT 732.970 0.010 733.970 4.280 ;
        RECT 734.810 0.010 735.810 4.280 ;
        RECT 736.650 0.010 737.650 4.280 ;
        RECT 738.490 0.010 739.490 4.280 ;
        RECT 740.330 0.010 741.330 4.280 ;
        RECT 742.170 0.010 743.170 4.280 ;
        RECT 744.010 0.010 745.010 4.280 ;
        RECT 745.850 0.010 746.850 4.280 ;
        RECT 747.690 0.010 748.690 4.280 ;
        RECT 749.530 0.010 750.530 4.280 ;
        RECT 751.370 0.010 752.370 4.280 ;
        RECT 753.210 0.010 754.210 4.280 ;
        RECT 755.050 0.010 756.050 4.280 ;
        RECT 756.890 0.010 757.890 4.280 ;
        RECT 758.730 0.010 759.730 4.280 ;
        RECT 760.570 0.010 761.570 4.280 ;
        RECT 762.410 0.010 763.410 4.280 ;
        RECT 764.250 0.010 765.250 4.280 ;
        RECT 766.090 0.010 767.090 4.280 ;
        RECT 767.930 0.010 768.930 4.280 ;
        RECT 769.770 0.010 770.770 4.280 ;
        RECT 771.610 0.010 772.610 4.280 ;
        RECT 773.450 0.010 774.450 4.280 ;
        RECT 775.290 0.010 776.290 4.280 ;
        RECT 777.130 0.010 778.130 4.280 ;
        RECT 778.970 0.010 779.970 4.280 ;
        RECT 780.810 0.010 781.350 4.280 ;
        RECT 782.190 0.010 783.190 4.280 ;
        RECT 784.030 0.010 785.030 4.280 ;
        RECT 785.870 0.010 786.870 4.280 ;
        RECT 787.710 0.010 788.710 4.280 ;
        RECT 789.550 0.010 790.550 4.280 ;
        RECT 791.390 0.010 792.390 4.280 ;
        RECT 793.230 0.010 794.230 4.280 ;
        RECT 795.070 0.010 796.070 4.280 ;
        RECT 796.910 0.010 797.910 4.280 ;
        RECT 798.750 0.010 799.750 4.280 ;
        RECT 800.590 0.010 801.590 4.280 ;
        RECT 802.430 0.010 803.430 4.280 ;
        RECT 804.270 0.010 805.270 4.280 ;
        RECT 806.110 0.010 807.110 4.280 ;
        RECT 807.950 0.010 808.950 4.280 ;
        RECT 809.790 0.010 810.790 4.280 ;
        RECT 811.630 0.010 812.630 4.280 ;
        RECT 813.470 0.010 814.470 4.280 ;
        RECT 815.310 0.010 816.310 4.280 ;
        RECT 817.150 0.010 818.150 4.280 ;
        RECT 818.990 0.010 819.990 4.280 ;
        RECT 820.830 0.010 821.830 4.280 ;
        RECT 822.670 0.010 823.670 4.280 ;
        RECT 824.510 0.010 825.510 4.280 ;
        RECT 826.350 0.010 827.350 4.280 ;
        RECT 828.190 0.010 829.190 4.280 ;
        RECT 830.030 0.010 831.030 4.280 ;
        RECT 831.870 0.010 832.870 4.280 ;
        RECT 833.710 0.010 834.710 4.280 ;
        RECT 835.550 0.010 836.550 4.280 ;
        RECT 837.390 0.010 838.390 4.280 ;
        RECT 839.230 0.010 840.230 4.280 ;
        RECT 841.070 0.010 841.610 4.280 ;
        RECT 842.450 0.010 843.450 4.280 ;
        RECT 844.290 0.010 845.290 4.280 ;
        RECT 846.130 0.010 847.130 4.280 ;
        RECT 847.970 0.010 848.970 4.280 ;
        RECT 849.810 0.010 850.810 4.280 ;
        RECT 851.650 0.010 852.650 4.280 ;
        RECT 853.490 0.010 854.490 4.280 ;
        RECT 855.330 0.010 856.330 4.280 ;
        RECT 857.170 0.010 858.170 4.280 ;
        RECT 859.010 0.010 860.010 4.280 ;
        RECT 860.850 0.010 861.850 4.280 ;
        RECT 862.690 0.010 863.690 4.280 ;
        RECT 864.530 0.010 865.530 4.280 ;
        RECT 866.370 0.010 867.370 4.280 ;
        RECT 868.210 0.010 869.210 4.280 ;
        RECT 870.050 0.010 871.050 4.280 ;
        RECT 871.890 0.010 872.890 4.280 ;
        RECT 873.730 0.010 874.730 4.280 ;
        RECT 875.570 0.010 876.570 4.280 ;
        RECT 877.410 0.010 878.410 4.280 ;
        RECT 879.250 0.010 880.250 4.280 ;
        RECT 881.090 0.010 882.090 4.280 ;
        RECT 882.930 0.010 883.930 4.280 ;
        RECT 884.770 0.010 885.770 4.280 ;
        RECT 886.610 0.010 887.610 4.280 ;
        RECT 888.450 0.010 889.450 4.280 ;
        RECT 890.290 0.010 891.290 4.280 ;
        RECT 892.130 0.010 893.130 4.280 ;
        RECT 893.970 0.010 894.970 4.280 ;
        RECT 895.810 0.010 896.810 4.280 ;
        RECT 897.650 0.010 898.650 4.280 ;
      LAYER met3 ;
        RECT 0.065 0.855 867.440 587.685 ;
      LAYER met4 ;
        RECT 239.495 10.240 251.040 265.705 ;
        RECT 253.440 10.240 327.840 265.705 ;
        RECT 330.240 10.240 404.640 265.705 ;
        RECT 407.040 10.240 479.025 265.705 ;
        RECT 239.495 0.855 479.025 10.240 ;
>>>>>>> 52a239652dd7a0722de75467858247e5f36b2500
  END
END user_proj_example
END LIBRARY

