magic
tech sky130A
magscale 1 2
timestamp 1623834721
<< obsli1 >>
rect 1104 1649 288880 287793
<< obsm1 >>
rect 290 688 289694 288040
<< metal2 >>
rect 1214 289200 1270 290000
rect 3698 289200 3754 290000
rect 6182 289200 6238 290000
rect 8666 289200 8722 290000
rect 11150 289200 11206 290000
rect 13634 289200 13690 290000
rect 16210 289200 16266 290000
rect 18694 289200 18750 290000
rect 21178 289200 21234 290000
rect 23662 289200 23718 290000
rect 26146 289200 26202 290000
rect 28630 289200 28686 290000
rect 31206 289200 31262 290000
rect 33690 289200 33746 290000
rect 36174 289200 36230 290000
rect 38658 289200 38714 290000
rect 41142 289200 41198 290000
rect 43626 289200 43682 290000
rect 46202 289200 46258 290000
rect 48686 289200 48742 290000
rect 51170 289200 51226 290000
rect 53654 289200 53710 290000
rect 56138 289200 56194 290000
rect 58622 289200 58678 290000
rect 61198 289200 61254 290000
rect 63682 289200 63738 290000
rect 66166 289200 66222 290000
rect 68650 289200 68706 290000
rect 71134 289200 71190 290000
rect 73710 289200 73766 290000
rect 76194 289200 76250 290000
rect 78678 289200 78734 290000
rect 81162 289200 81218 290000
rect 83646 289200 83702 290000
rect 86130 289200 86186 290000
rect 88706 289200 88762 290000
rect 91190 289200 91246 290000
rect 93674 289200 93730 290000
rect 96158 289200 96214 290000
rect 98642 289200 98698 290000
rect 101126 289200 101182 290000
rect 103702 289200 103758 290000
rect 106186 289200 106242 290000
rect 108670 289200 108726 290000
rect 111154 289200 111210 290000
rect 113638 289200 113694 290000
rect 116122 289200 116178 290000
rect 118698 289200 118754 290000
rect 121182 289200 121238 290000
rect 123666 289200 123722 290000
rect 126150 289200 126206 290000
rect 128634 289200 128690 290000
rect 131118 289200 131174 290000
rect 133694 289200 133750 290000
rect 136178 289200 136234 290000
rect 138662 289200 138718 290000
rect 141146 289200 141202 290000
rect 143630 289200 143686 290000
rect 146206 289200 146262 290000
rect 148690 289200 148746 290000
rect 151174 289200 151230 290000
rect 153658 289200 153714 290000
rect 156142 289200 156198 290000
rect 158626 289200 158682 290000
rect 161202 289200 161258 290000
rect 163686 289200 163742 290000
rect 166170 289200 166226 290000
rect 168654 289200 168710 290000
rect 171138 289200 171194 290000
rect 173622 289200 173678 290000
rect 176198 289200 176254 290000
rect 178682 289200 178738 290000
rect 181166 289200 181222 290000
rect 183650 289200 183706 290000
rect 186134 289200 186190 290000
rect 188618 289200 188674 290000
rect 191194 289200 191250 290000
rect 193678 289200 193734 290000
rect 196162 289200 196218 290000
rect 198646 289200 198702 290000
rect 201130 289200 201186 290000
rect 203614 289200 203670 290000
rect 206190 289200 206246 290000
rect 208674 289200 208730 290000
rect 211158 289200 211214 290000
rect 213642 289200 213698 290000
rect 216126 289200 216182 290000
rect 218702 289200 218758 290000
rect 221186 289200 221242 290000
rect 223670 289200 223726 290000
rect 226154 289200 226210 290000
rect 228638 289200 228694 290000
rect 231122 289200 231178 290000
rect 233698 289200 233754 290000
rect 236182 289200 236238 290000
rect 238666 289200 238722 290000
rect 241150 289200 241206 290000
rect 243634 289200 243690 290000
rect 246118 289200 246174 290000
rect 248694 289200 248750 290000
rect 251178 289200 251234 290000
rect 253662 289200 253718 290000
rect 256146 289200 256202 290000
rect 258630 289200 258686 290000
rect 261114 289200 261170 290000
rect 263690 289200 263746 290000
rect 266174 289200 266230 290000
rect 268658 289200 268714 290000
rect 271142 289200 271198 290000
rect 273626 289200 273682 290000
rect 276110 289200 276166 290000
rect 278686 289200 278742 290000
rect 281170 289200 281226 290000
rect 283654 289200 283710 290000
rect 286138 289200 286194 290000
rect 288622 289200 288678 290000
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 2042 0 2098 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3790 0 3846 800
rect 4434 0 4490 800
rect 4986 0 5042 800
rect 5538 0 5594 800
rect 6182 0 6238 800
rect 6734 0 6790 800
rect 7378 0 7434 800
rect 7930 0 7986 800
rect 8574 0 8630 800
rect 9126 0 9182 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11518 0 11574 800
rect 12070 0 12126 800
rect 12714 0 12770 800
rect 13266 0 13322 800
rect 13818 0 13874 800
rect 14462 0 14518 800
rect 15014 0 15070 800
rect 15658 0 15714 800
rect 16210 0 16266 800
rect 16854 0 16910 800
rect 17406 0 17462 800
rect 17958 0 18014 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19798 0 19854 800
rect 20350 0 20406 800
rect 20994 0 21050 800
rect 21546 0 21602 800
rect 22190 0 22246 800
rect 22742 0 22798 800
rect 23294 0 23350 800
rect 23938 0 23994 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25686 0 25742 800
rect 26330 0 26386 800
rect 26882 0 26938 800
rect 27434 0 27490 800
rect 28078 0 28134 800
rect 28630 0 28686 800
rect 29274 0 29330 800
rect 29826 0 29882 800
rect 30470 0 30526 800
rect 31022 0 31078 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32770 0 32826 800
rect 33414 0 33470 800
rect 33966 0 34022 800
rect 34610 0 34666 800
rect 35162 0 35218 800
rect 35714 0 35770 800
rect 36358 0 36414 800
rect 36910 0 36966 800
rect 37554 0 37610 800
rect 38106 0 38162 800
rect 38750 0 38806 800
rect 39302 0 39358 800
rect 39854 0 39910 800
rect 40498 0 40554 800
rect 41050 0 41106 800
rect 41694 0 41750 800
rect 42246 0 42302 800
rect 42890 0 42946 800
rect 43442 0 43498 800
rect 44086 0 44142 800
rect 44638 0 44694 800
rect 45190 0 45246 800
rect 45834 0 45890 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 47582 0 47638 800
rect 48226 0 48282 800
rect 48778 0 48834 800
rect 49330 0 49386 800
rect 49974 0 50030 800
rect 50526 0 50582 800
rect 51170 0 51226 800
rect 51722 0 51778 800
rect 52366 0 52422 800
rect 52918 0 52974 800
rect 53470 0 53526 800
rect 54114 0 54170 800
rect 54666 0 54722 800
rect 55310 0 55366 800
rect 55862 0 55918 800
rect 56506 0 56562 800
rect 57058 0 57114 800
rect 57610 0 57666 800
rect 58254 0 58310 800
rect 58806 0 58862 800
rect 59450 0 59506 800
rect 60002 0 60058 800
rect 60646 0 60702 800
rect 61198 0 61254 800
rect 61750 0 61806 800
rect 62394 0 62450 800
rect 62946 0 63002 800
rect 63590 0 63646 800
rect 64142 0 64198 800
rect 64786 0 64842 800
rect 65338 0 65394 800
rect 65982 0 66038 800
rect 66534 0 66590 800
rect 67086 0 67142 800
rect 67730 0 67786 800
rect 68282 0 68338 800
rect 68926 0 68982 800
rect 69478 0 69534 800
rect 70122 0 70178 800
rect 70674 0 70730 800
rect 71226 0 71282 800
rect 71870 0 71926 800
rect 72422 0 72478 800
rect 73066 0 73122 800
rect 73618 0 73674 800
rect 74262 0 74318 800
rect 74814 0 74870 800
rect 75366 0 75422 800
rect 76010 0 76066 800
rect 76562 0 76618 800
rect 77206 0 77262 800
rect 77758 0 77814 800
rect 78402 0 78458 800
rect 78954 0 79010 800
rect 79506 0 79562 800
rect 80150 0 80206 800
rect 80702 0 80758 800
rect 81346 0 81402 800
rect 81898 0 81954 800
rect 82542 0 82598 800
rect 83094 0 83150 800
rect 83738 0 83794 800
rect 84290 0 84346 800
rect 84842 0 84898 800
rect 85486 0 85542 800
rect 86038 0 86094 800
rect 86682 0 86738 800
rect 87234 0 87290 800
rect 87878 0 87934 800
rect 88430 0 88486 800
rect 88982 0 89038 800
rect 89626 0 89682 800
rect 90178 0 90234 800
rect 90822 0 90878 800
rect 91374 0 91430 800
rect 92018 0 92074 800
rect 92570 0 92626 800
rect 93122 0 93178 800
rect 93766 0 93822 800
rect 94318 0 94374 800
rect 94962 0 95018 800
rect 95514 0 95570 800
rect 96158 0 96214 800
rect 96710 0 96766 800
rect 97262 0 97318 800
rect 97906 0 97962 800
rect 98458 0 98514 800
rect 99102 0 99158 800
rect 99654 0 99710 800
rect 100298 0 100354 800
rect 100850 0 100906 800
rect 101402 0 101458 800
rect 102046 0 102102 800
rect 102598 0 102654 800
rect 103242 0 103298 800
rect 103794 0 103850 800
rect 104438 0 104494 800
rect 104990 0 105046 800
rect 105634 0 105690 800
rect 106186 0 106242 800
rect 106738 0 106794 800
rect 107382 0 107438 800
rect 107934 0 107990 800
rect 108578 0 108634 800
rect 109130 0 109186 800
rect 109774 0 109830 800
rect 110326 0 110382 800
rect 110878 0 110934 800
rect 111522 0 111578 800
rect 112074 0 112130 800
rect 112718 0 112774 800
rect 113270 0 113326 800
rect 113914 0 113970 800
rect 114466 0 114522 800
rect 115018 0 115074 800
rect 115662 0 115718 800
rect 116214 0 116270 800
rect 116858 0 116914 800
rect 117410 0 117466 800
rect 118054 0 118110 800
rect 118606 0 118662 800
rect 119158 0 119214 800
rect 119802 0 119858 800
rect 120354 0 120410 800
rect 120998 0 121054 800
rect 121550 0 121606 800
rect 122194 0 122250 800
rect 122746 0 122802 800
rect 123298 0 123354 800
rect 123942 0 123998 800
rect 124494 0 124550 800
rect 125138 0 125194 800
rect 125690 0 125746 800
rect 126334 0 126390 800
rect 126886 0 126942 800
rect 127530 0 127586 800
rect 128082 0 128138 800
rect 128634 0 128690 800
rect 129278 0 129334 800
rect 129830 0 129886 800
rect 130474 0 130530 800
rect 131026 0 131082 800
rect 131670 0 131726 800
rect 132222 0 132278 800
rect 132774 0 132830 800
rect 133418 0 133474 800
rect 133970 0 134026 800
rect 134614 0 134670 800
rect 135166 0 135222 800
rect 135810 0 135866 800
rect 136362 0 136418 800
rect 136914 0 136970 800
rect 137558 0 137614 800
rect 138110 0 138166 800
rect 138754 0 138810 800
rect 139306 0 139362 800
rect 139950 0 140006 800
rect 140502 0 140558 800
rect 141054 0 141110 800
rect 141698 0 141754 800
rect 142250 0 142306 800
rect 142894 0 142950 800
rect 143446 0 143502 800
rect 144090 0 144146 800
rect 144642 0 144698 800
rect 145286 0 145342 800
rect 145838 0 145894 800
rect 146390 0 146446 800
rect 147034 0 147090 800
rect 147586 0 147642 800
rect 148230 0 148286 800
rect 148782 0 148838 800
rect 149426 0 149482 800
rect 149978 0 150034 800
rect 150530 0 150586 800
rect 151174 0 151230 800
rect 151726 0 151782 800
rect 152370 0 152426 800
rect 152922 0 152978 800
rect 153566 0 153622 800
rect 154118 0 154174 800
rect 154670 0 154726 800
rect 155314 0 155370 800
rect 155866 0 155922 800
rect 156510 0 156566 800
rect 157062 0 157118 800
rect 157706 0 157762 800
rect 158258 0 158314 800
rect 158810 0 158866 800
rect 159454 0 159510 800
rect 160006 0 160062 800
rect 160650 0 160706 800
rect 161202 0 161258 800
rect 161846 0 161902 800
rect 162398 0 162454 800
rect 162950 0 163006 800
rect 163594 0 163650 800
rect 164146 0 164202 800
rect 164790 0 164846 800
rect 165342 0 165398 800
rect 165986 0 166042 800
rect 166538 0 166594 800
rect 167182 0 167238 800
rect 167734 0 167790 800
rect 168286 0 168342 800
rect 168930 0 168986 800
rect 169482 0 169538 800
rect 170126 0 170182 800
rect 170678 0 170734 800
rect 171322 0 171378 800
rect 171874 0 171930 800
rect 172426 0 172482 800
rect 173070 0 173126 800
rect 173622 0 173678 800
rect 174266 0 174322 800
rect 174818 0 174874 800
rect 175462 0 175518 800
rect 176014 0 176070 800
rect 176566 0 176622 800
rect 177210 0 177266 800
rect 177762 0 177818 800
rect 178406 0 178462 800
rect 178958 0 179014 800
rect 179602 0 179658 800
rect 180154 0 180210 800
rect 180706 0 180762 800
rect 181350 0 181406 800
rect 181902 0 181958 800
rect 182546 0 182602 800
rect 183098 0 183154 800
rect 183742 0 183798 800
rect 184294 0 184350 800
rect 184846 0 184902 800
rect 185490 0 185546 800
rect 186042 0 186098 800
rect 186686 0 186742 800
rect 187238 0 187294 800
rect 187882 0 187938 800
rect 188434 0 188490 800
rect 189078 0 189134 800
rect 189630 0 189686 800
rect 190182 0 190238 800
rect 190826 0 190882 800
rect 191378 0 191434 800
rect 192022 0 192078 800
rect 192574 0 192630 800
rect 193218 0 193274 800
rect 193770 0 193826 800
rect 194322 0 194378 800
rect 194966 0 195022 800
rect 195518 0 195574 800
rect 196162 0 196218 800
rect 196714 0 196770 800
rect 197358 0 197414 800
rect 197910 0 197966 800
rect 198462 0 198518 800
rect 199106 0 199162 800
rect 199658 0 199714 800
rect 200302 0 200358 800
rect 200854 0 200910 800
rect 201498 0 201554 800
rect 202050 0 202106 800
rect 202602 0 202658 800
rect 203246 0 203302 800
rect 203798 0 203854 800
rect 204442 0 204498 800
rect 204994 0 205050 800
rect 205638 0 205694 800
rect 206190 0 206246 800
rect 206742 0 206798 800
rect 207386 0 207442 800
rect 207938 0 207994 800
rect 208582 0 208638 800
rect 209134 0 209190 800
rect 209778 0 209834 800
rect 210330 0 210386 800
rect 210974 0 211030 800
rect 211526 0 211582 800
rect 212078 0 212134 800
rect 212722 0 212778 800
rect 213274 0 213330 800
rect 213918 0 213974 800
rect 214470 0 214526 800
rect 215114 0 215170 800
rect 215666 0 215722 800
rect 216218 0 216274 800
rect 216862 0 216918 800
rect 217414 0 217470 800
rect 218058 0 218114 800
rect 218610 0 218666 800
rect 219254 0 219310 800
rect 219806 0 219862 800
rect 220358 0 220414 800
rect 221002 0 221058 800
rect 221554 0 221610 800
rect 222198 0 222254 800
rect 222750 0 222806 800
rect 223394 0 223450 800
rect 223946 0 224002 800
rect 224498 0 224554 800
rect 225142 0 225198 800
rect 225694 0 225750 800
rect 226338 0 226394 800
rect 226890 0 226946 800
rect 227534 0 227590 800
rect 228086 0 228142 800
rect 228730 0 228786 800
rect 229282 0 229338 800
rect 229834 0 229890 800
rect 230478 0 230534 800
rect 231030 0 231086 800
rect 231674 0 231730 800
rect 232226 0 232282 800
rect 232870 0 232926 800
rect 233422 0 233478 800
rect 233974 0 234030 800
rect 234618 0 234674 800
rect 235170 0 235226 800
rect 235814 0 235870 800
rect 236366 0 236422 800
rect 237010 0 237066 800
rect 237562 0 237618 800
rect 238114 0 238170 800
rect 238758 0 238814 800
rect 239310 0 239366 800
rect 239954 0 240010 800
rect 240506 0 240562 800
rect 241150 0 241206 800
rect 241702 0 241758 800
rect 242254 0 242310 800
rect 242898 0 242954 800
rect 243450 0 243506 800
rect 244094 0 244150 800
rect 244646 0 244702 800
rect 245290 0 245346 800
rect 245842 0 245898 800
rect 246394 0 246450 800
rect 247038 0 247094 800
rect 247590 0 247646 800
rect 248234 0 248290 800
rect 248786 0 248842 800
rect 249430 0 249486 800
rect 249982 0 250038 800
rect 250626 0 250682 800
rect 251178 0 251234 800
rect 251730 0 251786 800
rect 252374 0 252430 800
rect 252926 0 252982 800
rect 253570 0 253626 800
rect 254122 0 254178 800
rect 254766 0 254822 800
rect 255318 0 255374 800
rect 255870 0 255926 800
rect 256514 0 256570 800
rect 257066 0 257122 800
rect 257710 0 257766 800
rect 258262 0 258318 800
rect 258906 0 258962 800
rect 259458 0 259514 800
rect 260010 0 260066 800
rect 260654 0 260710 800
rect 261206 0 261262 800
rect 261850 0 261906 800
rect 262402 0 262458 800
rect 263046 0 263102 800
rect 263598 0 263654 800
rect 264150 0 264206 800
rect 264794 0 264850 800
rect 265346 0 265402 800
rect 265990 0 266046 800
rect 266542 0 266598 800
rect 267186 0 267242 800
rect 267738 0 267794 800
rect 268290 0 268346 800
rect 268934 0 268990 800
rect 269486 0 269542 800
rect 270130 0 270186 800
rect 270682 0 270738 800
rect 271326 0 271382 800
rect 271878 0 271934 800
rect 272522 0 272578 800
rect 273074 0 273130 800
rect 273626 0 273682 800
rect 274270 0 274326 800
rect 274822 0 274878 800
rect 275466 0 275522 800
rect 276018 0 276074 800
rect 276662 0 276718 800
rect 277214 0 277270 800
rect 277766 0 277822 800
rect 278410 0 278466 800
rect 278962 0 279018 800
rect 279606 0 279662 800
rect 280158 0 280214 800
rect 280802 0 280858 800
rect 281354 0 281410 800
rect 281906 0 281962 800
rect 282550 0 282606 800
rect 283102 0 283158 800
rect 283746 0 283802 800
rect 284298 0 284354 800
rect 284942 0 284998 800
rect 285494 0 285550 800
rect 286046 0 286102 800
rect 286690 0 286746 800
rect 287242 0 287298 800
rect 287886 0 287942 800
rect 288438 0 288494 800
rect 289082 0 289138 800
rect 289634 0 289690 800
<< obsm2 >>
rect 296 289144 1158 289200
rect 1326 289144 3642 289200
rect 3810 289144 6126 289200
rect 6294 289144 8610 289200
rect 8778 289144 11094 289200
rect 11262 289144 13578 289200
rect 13746 289144 16154 289200
rect 16322 289144 18638 289200
rect 18806 289144 21122 289200
rect 21290 289144 23606 289200
rect 23774 289144 26090 289200
rect 26258 289144 28574 289200
rect 28742 289144 31150 289200
rect 31318 289144 33634 289200
rect 33802 289144 36118 289200
rect 36286 289144 38602 289200
rect 38770 289144 41086 289200
rect 41254 289144 43570 289200
rect 43738 289144 46146 289200
rect 46314 289144 48630 289200
rect 48798 289144 51114 289200
rect 51282 289144 53598 289200
rect 53766 289144 56082 289200
rect 56250 289144 58566 289200
rect 58734 289144 61142 289200
rect 61310 289144 63626 289200
rect 63794 289144 66110 289200
rect 66278 289144 68594 289200
rect 68762 289144 71078 289200
rect 71246 289144 73654 289200
rect 73822 289144 76138 289200
rect 76306 289144 78622 289200
rect 78790 289144 81106 289200
rect 81274 289144 83590 289200
rect 83758 289144 86074 289200
rect 86242 289144 88650 289200
rect 88818 289144 91134 289200
rect 91302 289144 93618 289200
rect 93786 289144 96102 289200
rect 96270 289144 98586 289200
rect 98754 289144 101070 289200
rect 101238 289144 103646 289200
rect 103814 289144 106130 289200
rect 106298 289144 108614 289200
rect 108782 289144 111098 289200
rect 111266 289144 113582 289200
rect 113750 289144 116066 289200
rect 116234 289144 118642 289200
rect 118810 289144 121126 289200
rect 121294 289144 123610 289200
rect 123778 289144 126094 289200
rect 126262 289144 128578 289200
rect 128746 289144 131062 289200
rect 131230 289144 133638 289200
rect 133806 289144 136122 289200
rect 136290 289144 138606 289200
rect 138774 289144 141090 289200
rect 141258 289144 143574 289200
rect 143742 289144 146150 289200
rect 146318 289144 148634 289200
rect 148802 289144 151118 289200
rect 151286 289144 153602 289200
rect 153770 289144 156086 289200
rect 156254 289144 158570 289200
rect 158738 289144 161146 289200
rect 161314 289144 163630 289200
rect 163798 289144 166114 289200
rect 166282 289144 168598 289200
rect 168766 289144 171082 289200
rect 171250 289144 173566 289200
rect 173734 289144 176142 289200
rect 176310 289144 178626 289200
rect 178794 289144 181110 289200
rect 181278 289144 183594 289200
rect 183762 289144 186078 289200
rect 186246 289144 188562 289200
rect 188730 289144 191138 289200
rect 191306 289144 193622 289200
rect 193790 289144 196106 289200
rect 196274 289144 198590 289200
rect 198758 289144 201074 289200
rect 201242 289144 203558 289200
rect 203726 289144 206134 289200
rect 206302 289144 208618 289200
rect 208786 289144 211102 289200
rect 211270 289144 213586 289200
rect 213754 289144 216070 289200
rect 216238 289144 218646 289200
rect 218814 289144 221130 289200
rect 221298 289144 223614 289200
rect 223782 289144 226098 289200
rect 226266 289144 228582 289200
rect 228750 289144 231066 289200
rect 231234 289144 233642 289200
rect 233810 289144 236126 289200
rect 236294 289144 238610 289200
rect 238778 289144 241094 289200
rect 241262 289144 243578 289200
rect 243746 289144 246062 289200
rect 246230 289144 248638 289200
rect 248806 289144 251122 289200
rect 251290 289144 253606 289200
rect 253774 289144 256090 289200
rect 256258 289144 258574 289200
rect 258742 289144 261058 289200
rect 261226 289144 263634 289200
rect 263802 289144 266118 289200
rect 266286 289144 268602 289200
rect 268770 289144 271086 289200
rect 271254 289144 273570 289200
rect 273738 289144 276054 289200
rect 276222 289144 278630 289200
rect 278798 289144 281114 289200
rect 281282 289144 283598 289200
rect 283766 289144 286082 289200
rect 286250 289144 288566 289200
rect 288734 289144 289688 289200
rect 296 856 289688 289144
rect 406 682 790 856
rect 958 682 1342 856
rect 1510 682 1986 856
rect 2154 682 2538 856
rect 2706 682 3182 856
rect 3350 682 3734 856
rect 3902 682 4378 856
rect 4546 682 4930 856
rect 5098 682 5482 856
rect 5650 682 6126 856
rect 6294 682 6678 856
rect 6846 682 7322 856
rect 7490 682 7874 856
rect 8042 682 8518 856
rect 8686 682 9070 856
rect 9238 682 9622 856
rect 9790 682 10266 856
rect 10434 682 10818 856
rect 10986 682 11462 856
rect 11630 682 12014 856
rect 12182 682 12658 856
rect 12826 682 13210 856
rect 13378 682 13762 856
rect 13930 682 14406 856
rect 14574 682 14958 856
rect 15126 682 15602 856
rect 15770 682 16154 856
rect 16322 682 16798 856
rect 16966 682 17350 856
rect 17518 682 17902 856
rect 18070 682 18546 856
rect 18714 682 19098 856
rect 19266 682 19742 856
rect 19910 682 20294 856
rect 20462 682 20938 856
rect 21106 682 21490 856
rect 21658 682 22134 856
rect 22302 682 22686 856
rect 22854 682 23238 856
rect 23406 682 23882 856
rect 24050 682 24434 856
rect 24602 682 25078 856
rect 25246 682 25630 856
rect 25798 682 26274 856
rect 26442 682 26826 856
rect 26994 682 27378 856
rect 27546 682 28022 856
rect 28190 682 28574 856
rect 28742 682 29218 856
rect 29386 682 29770 856
rect 29938 682 30414 856
rect 30582 682 30966 856
rect 31134 682 31518 856
rect 31686 682 32162 856
rect 32330 682 32714 856
rect 32882 682 33358 856
rect 33526 682 33910 856
rect 34078 682 34554 856
rect 34722 682 35106 856
rect 35274 682 35658 856
rect 35826 682 36302 856
rect 36470 682 36854 856
rect 37022 682 37498 856
rect 37666 682 38050 856
rect 38218 682 38694 856
rect 38862 682 39246 856
rect 39414 682 39798 856
rect 39966 682 40442 856
rect 40610 682 40994 856
rect 41162 682 41638 856
rect 41806 682 42190 856
rect 42358 682 42834 856
rect 43002 682 43386 856
rect 43554 682 44030 856
rect 44198 682 44582 856
rect 44750 682 45134 856
rect 45302 682 45778 856
rect 45946 682 46330 856
rect 46498 682 46974 856
rect 47142 682 47526 856
rect 47694 682 48170 856
rect 48338 682 48722 856
rect 48890 682 49274 856
rect 49442 682 49918 856
rect 50086 682 50470 856
rect 50638 682 51114 856
rect 51282 682 51666 856
rect 51834 682 52310 856
rect 52478 682 52862 856
rect 53030 682 53414 856
rect 53582 682 54058 856
rect 54226 682 54610 856
rect 54778 682 55254 856
rect 55422 682 55806 856
rect 55974 682 56450 856
rect 56618 682 57002 856
rect 57170 682 57554 856
rect 57722 682 58198 856
rect 58366 682 58750 856
rect 58918 682 59394 856
rect 59562 682 59946 856
rect 60114 682 60590 856
rect 60758 682 61142 856
rect 61310 682 61694 856
rect 61862 682 62338 856
rect 62506 682 62890 856
rect 63058 682 63534 856
rect 63702 682 64086 856
rect 64254 682 64730 856
rect 64898 682 65282 856
rect 65450 682 65926 856
rect 66094 682 66478 856
rect 66646 682 67030 856
rect 67198 682 67674 856
rect 67842 682 68226 856
rect 68394 682 68870 856
rect 69038 682 69422 856
rect 69590 682 70066 856
rect 70234 682 70618 856
rect 70786 682 71170 856
rect 71338 682 71814 856
rect 71982 682 72366 856
rect 72534 682 73010 856
rect 73178 682 73562 856
rect 73730 682 74206 856
rect 74374 682 74758 856
rect 74926 682 75310 856
rect 75478 682 75954 856
rect 76122 682 76506 856
rect 76674 682 77150 856
rect 77318 682 77702 856
rect 77870 682 78346 856
rect 78514 682 78898 856
rect 79066 682 79450 856
rect 79618 682 80094 856
rect 80262 682 80646 856
rect 80814 682 81290 856
rect 81458 682 81842 856
rect 82010 682 82486 856
rect 82654 682 83038 856
rect 83206 682 83682 856
rect 83850 682 84234 856
rect 84402 682 84786 856
rect 84954 682 85430 856
rect 85598 682 85982 856
rect 86150 682 86626 856
rect 86794 682 87178 856
rect 87346 682 87822 856
rect 87990 682 88374 856
rect 88542 682 88926 856
rect 89094 682 89570 856
rect 89738 682 90122 856
rect 90290 682 90766 856
rect 90934 682 91318 856
rect 91486 682 91962 856
rect 92130 682 92514 856
rect 92682 682 93066 856
rect 93234 682 93710 856
rect 93878 682 94262 856
rect 94430 682 94906 856
rect 95074 682 95458 856
rect 95626 682 96102 856
rect 96270 682 96654 856
rect 96822 682 97206 856
rect 97374 682 97850 856
rect 98018 682 98402 856
rect 98570 682 99046 856
rect 99214 682 99598 856
rect 99766 682 100242 856
rect 100410 682 100794 856
rect 100962 682 101346 856
rect 101514 682 101990 856
rect 102158 682 102542 856
rect 102710 682 103186 856
rect 103354 682 103738 856
rect 103906 682 104382 856
rect 104550 682 104934 856
rect 105102 682 105578 856
rect 105746 682 106130 856
rect 106298 682 106682 856
rect 106850 682 107326 856
rect 107494 682 107878 856
rect 108046 682 108522 856
rect 108690 682 109074 856
rect 109242 682 109718 856
rect 109886 682 110270 856
rect 110438 682 110822 856
rect 110990 682 111466 856
rect 111634 682 112018 856
rect 112186 682 112662 856
rect 112830 682 113214 856
rect 113382 682 113858 856
rect 114026 682 114410 856
rect 114578 682 114962 856
rect 115130 682 115606 856
rect 115774 682 116158 856
rect 116326 682 116802 856
rect 116970 682 117354 856
rect 117522 682 117998 856
rect 118166 682 118550 856
rect 118718 682 119102 856
rect 119270 682 119746 856
rect 119914 682 120298 856
rect 120466 682 120942 856
rect 121110 682 121494 856
rect 121662 682 122138 856
rect 122306 682 122690 856
rect 122858 682 123242 856
rect 123410 682 123886 856
rect 124054 682 124438 856
rect 124606 682 125082 856
rect 125250 682 125634 856
rect 125802 682 126278 856
rect 126446 682 126830 856
rect 126998 682 127474 856
rect 127642 682 128026 856
rect 128194 682 128578 856
rect 128746 682 129222 856
rect 129390 682 129774 856
rect 129942 682 130418 856
rect 130586 682 130970 856
rect 131138 682 131614 856
rect 131782 682 132166 856
rect 132334 682 132718 856
rect 132886 682 133362 856
rect 133530 682 133914 856
rect 134082 682 134558 856
rect 134726 682 135110 856
rect 135278 682 135754 856
rect 135922 682 136306 856
rect 136474 682 136858 856
rect 137026 682 137502 856
rect 137670 682 138054 856
rect 138222 682 138698 856
rect 138866 682 139250 856
rect 139418 682 139894 856
rect 140062 682 140446 856
rect 140614 682 140998 856
rect 141166 682 141642 856
rect 141810 682 142194 856
rect 142362 682 142838 856
rect 143006 682 143390 856
rect 143558 682 144034 856
rect 144202 682 144586 856
rect 144754 682 145230 856
rect 145398 682 145782 856
rect 145950 682 146334 856
rect 146502 682 146978 856
rect 147146 682 147530 856
rect 147698 682 148174 856
rect 148342 682 148726 856
rect 148894 682 149370 856
rect 149538 682 149922 856
rect 150090 682 150474 856
rect 150642 682 151118 856
rect 151286 682 151670 856
rect 151838 682 152314 856
rect 152482 682 152866 856
rect 153034 682 153510 856
rect 153678 682 154062 856
rect 154230 682 154614 856
rect 154782 682 155258 856
rect 155426 682 155810 856
rect 155978 682 156454 856
rect 156622 682 157006 856
rect 157174 682 157650 856
rect 157818 682 158202 856
rect 158370 682 158754 856
rect 158922 682 159398 856
rect 159566 682 159950 856
rect 160118 682 160594 856
rect 160762 682 161146 856
rect 161314 682 161790 856
rect 161958 682 162342 856
rect 162510 682 162894 856
rect 163062 682 163538 856
rect 163706 682 164090 856
rect 164258 682 164734 856
rect 164902 682 165286 856
rect 165454 682 165930 856
rect 166098 682 166482 856
rect 166650 682 167126 856
rect 167294 682 167678 856
rect 167846 682 168230 856
rect 168398 682 168874 856
rect 169042 682 169426 856
rect 169594 682 170070 856
rect 170238 682 170622 856
rect 170790 682 171266 856
rect 171434 682 171818 856
rect 171986 682 172370 856
rect 172538 682 173014 856
rect 173182 682 173566 856
rect 173734 682 174210 856
rect 174378 682 174762 856
rect 174930 682 175406 856
rect 175574 682 175958 856
rect 176126 682 176510 856
rect 176678 682 177154 856
rect 177322 682 177706 856
rect 177874 682 178350 856
rect 178518 682 178902 856
rect 179070 682 179546 856
rect 179714 682 180098 856
rect 180266 682 180650 856
rect 180818 682 181294 856
rect 181462 682 181846 856
rect 182014 682 182490 856
rect 182658 682 183042 856
rect 183210 682 183686 856
rect 183854 682 184238 856
rect 184406 682 184790 856
rect 184958 682 185434 856
rect 185602 682 185986 856
rect 186154 682 186630 856
rect 186798 682 187182 856
rect 187350 682 187826 856
rect 187994 682 188378 856
rect 188546 682 189022 856
rect 189190 682 189574 856
rect 189742 682 190126 856
rect 190294 682 190770 856
rect 190938 682 191322 856
rect 191490 682 191966 856
rect 192134 682 192518 856
rect 192686 682 193162 856
rect 193330 682 193714 856
rect 193882 682 194266 856
rect 194434 682 194910 856
rect 195078 682 195462 856
rect 195630 682 196106 856
rect 196274 682 196658 856
rect 196826 682 197302 856
rect 197470 682 197854 856
rect 198022 682 198406 856
rect 198574 682 199050 856
rect 199218 682 199602 856
rect 199770 682 200246 856
rect 200414 682 200798 856
rect 200966 682 201442 856
rect 201610 682 201994 856
rect 202162 682 202546 856
rect 202714 682 203190 856
rect 203358 682 203742 856
rect 203910 682 204386 856
rect 204554 682 204938 856
rect 205106 682 205582 856
rect 205750 682 206134 856
rect 206302 682 206686 856
rect 206854 682 207330 856
rect 207498 682 207882 856
rect 208050 682 208526 856
rect 208694 682 209078 856
rect 209246 682 209722 856
rect 209890 682 210274 856
rect 210442 682 210918 856
rect 211086 682 211470 856
rect 211638 682 212022 856
rect 212190 682 212666 856
rect 212834 682 213218 856
rect 213386 682 213862 856
rect 214030 682 214414 856
rect 214582 682 215058 856
rect 215226 682 215610 856
rect 215778 682 216162 856
rect 216330 682 216806 856
rect 216974 682 217358 856
rect 217526 682 218002 856
rect 218170 682 218554 856
rect 218722 682 219198 856
rect 219366 682 219750 856
rect 219918 682 220302 856
rect 220470 682 220946 856
rect 221114 682 221498 856
rect 221666 682 222142 856
rect 222310 682 222694 856
rect 222862 682 223338 856
rect 223506 682 223890 856
rect 224058 682 224442 856
rect 224610 682 225086 856
rect 225254 682 225638 856
rect 225806 682 226282 856
rect 226450 682 226834 856
rect 227002 682 227478 856
rect 227646 682 228030 856
rect 228198 682 228674 856
rect 228842 682 229226 856
rect 229394 682 229778 856
rect 229946 682 230422 856
rect 230590 682 230974 856
rect 231142 682 231618 856
rect 231786 682 232170 856
rect 232338 682 232814 856
rect 232982 682 233366 856
rect 233534 682 233918 856
rect 234086 682 234562 856
rect 234730 682 235114 856
rect 235282 682 235758 856
rect 235926 682 236310 856
rect 236478 682 236954 856
rect 237122 682 237506 856
rect 237674 682 238058 856
rect 238226 682 238702 856
rect 238870 682 239254 856
rect 239422 682 239898 856
rect 240066 682 240450 856
rect 240618 682 241094 856
rect 241262 682 241646 856
rect 241814 682 242198 856
rect 242366 682 242842 856
rect 243010 682 243394 856
rect 243562 682 244038 856
rect 244206 682 244590 856
rect 244758 682 245234 856
rect 245402 682 245786 856
rect 245954 682 246338 856
rect 246506 682 246982 856
rect 247150 682 247534 856
rect 247702 682 248178 856
rect 248346 682 248730 856
rect 248898 682 249374 856
rect 249542 682 249926 856
rect 250094 682 250570 856
rect 250738 682 251122 856
rect 251290 682 251674 856
rect 251842 682 252318 856
rect 252486 682 252870 856
rect 253038 682 253514 856
rect 253682 682 254066 856
rect 254234 682 254710 856
rect 254878 682 255262 856
rect 255430 682 255814 856
rect 255982 682 256458 856
rect 256626 682 257010 856
rect 257178 682 257654 856
rect 257822 682 258206 856
rect 258374 682 258850 856
rect 259018 682 259402 856
rect 259570 682 259954 856
rect 260122 682 260598 856
rect 260766 682 261150 856
rect 261318 682 261794 856
rect 261962 682 262346 856
rect 262514 682 262990 856
rect 263158 682 263542 856
rect 263710 682 264094 856
rect 264262 682 264738 856
rect 264906 682 265290 856
rect 265458 682 265934 856
rect 266102 682 266486 856
rect 266654 682 267130 856
rect 267298 682 267682 856
rect 267850 682 268234 856
rect 268402 682 268878 856
rect 269046 682 269430 856
rect 269598 682 270074 856
rect 270242 682 270626 856
rect 270794 682 271270 856
rect 271438 682 271822 856
rect 271990 682 272466 856
rect 272634 682 273018 856
rect 273186 682 273570 856
rect 273738 682 274214 856
rect 274382 682 274766 856
rect 274934 682 275410 856
rect 275578 682 275962 856
rect 276130 682 276606 856
rect 276774 682 277158 856
rect 277326 682 277710 856
rect 277878 682 278354 856
rect 278522 682 278906 856
rect 279074 682 279550 856
rect 279718 682 280102 856
rect 280270 682 280746 856
rect 280914 682 281298 856
rect 281466 682 281850 856
rect 282018 682 282494 856
rect 282662 682 283046 856
rect 283214 682 283690 856
rect 283858 682 284242 856
rect 284410 682 284886 856
rect 285054 682 285438 856
rect 285606 682 285990 856
rect 286158 682 286634 856
rect 286802 682 287186 856
rect 287354 682 287830 856
rect 287998 682 288382 856
rect 288550 682 289026 856
rect 289194 682 289578 856
<< metal3 >>
rect 0 217472 800 217592
rect 0 72496 800 72616
<< obsm3 >>
rect 800 217672 288315 287809
rect 880 217392 288315 217672
rect 800 72696 288315 217392
rect 880 72416 288315 72696
rect 800 2143 288315 72416
<< metal4 >>
rect 4208 2128 4528 287824
rect 4868 2176 5188 287776
rect 5528 2176 5848 287776
rect 6188 2176 6508 287776
rect 19568 2128 19888 287824
rect 20228 2176 20548 287776
rect 20888 2176 21208 287776
rect 21548 2176 21868 287776
rect 34928 2128 35248 287824
rect 35588 2176 35908 287776
rect 36248 2176 36568 287776
rect 36908 2176 37228 287776
rect 50288 2128 50608 287824
rect 50948 2176 51268 287776
rect 51608 2176 51928 287776
rect 52268 2176 52588 287776
rect 65648 2128 65968 287824
rect 66308 2176 66628 287776
rect 66968 2176 67288 287776
rect 67628 2176 67948 287776
rect 81008 2128 81328 287824
rect 81668 2176 81988 287776
rect 82328 2176 82648 287776
rect 82988 2176 83308 287776
rect 96368 2128 96688 287824
rect 97028 2176 97348 287776
rect 97688 2176 98008 287776
rect 98348 2176 98668 287776
rect 111728 2128 112048 287824
rect 112388 2176 112708 287776
rect 113048 2176 113368 287776
rect 113708 2176 114028 287776
rect 127088 2128 127408 287824
rect 127748 2176 128068 287776
rect 128408 2176 128728 287776
rect 129068 2176 129388 287776
rect 142448 2128 142768 287824
rect 143108 2176 143428 287776
rect 143768 2176 144088 287776
rect 144428 2176 144748 287776
rect 157808 2128 158128 287824
rect 158468 2176 158788 287776
rect 159128 2176 159448 287776
rect 159788 2176 160108 287776
rect 173168 2128 173488 287824
rect 173828 2176 174148 287776
rect 174488 2176 174808 287776
rect 175148 2176 175468 287776
rect 188528 2128 188848 287824
rect 189188 2176 189508 287776
rect 189848 2176 190168 287776
rect 190508 2176 190828 287776
rect 203888 2128 204208 287824
rect 204548 2176 204868 287776
rect 205208 2176 205528 287776
rect 205868 2176 206188 287776
rect 219248 2128 219568 287824
rect 219908 2176 220228 287776
rect 220568 2176 220888 287776
rect 221228 2176 221548 287776
rect 234608 2128 234928 287824
rect 235268 2176 235588 287776
rect 235928 2176 236248 287776
rect 236588 2176 236908 287776
rect 249968 2128 250288 287824
rect 250628 2176 250948 287776
rect 251288 2176 251608 287776
rect 251948 2176 252268 287776
rect 265328 2128 265648 287824
rect 265988 2176 266308 287776
rect 266648 2176 266968 287776
rect 267308 2176 267628 287776
rect 280688 2128 281008 287824
rect 281348 2176 281668 287776
rect 282008 2176 282328 287776
rect 282668 2176 282988 287776
<< obsm4 >>
rect 9627 2619 19488 287605
rect 19968 2619 20148 287605
rect 20628 2619 20808 287605
rect 21288 2619 21468 287605
rect 21948 2619 34848 287605
rect 35328 2619 35508 287605
rect 35988 2619 36168 287605
rect 36648 2619 36828 287605
rect 37308 2619 50208 287605
rect 50688 2619 50868 287605
rect 51348 2619 51528 287605
rect 52008 2619 52188 287605
rect 52668 2619 65568 287605
rect 66048 2619 66228 287605
rect 66708 2619 66888 287605
rect 67368 2619 67548 287605
rect 68028 2619 80928 287605
rect 81408 2619 81588 287605
rect 82068 2619 82248 287605
rect 82728 2619 82908 287605
rect 83388 2619 96288 287605
rect 96768 2619 96948 287605
rect 97428 2619 97608 287605
rect 98088 2619 98268 287605
rect 98748 2619 111648 287605
rect 112128 2619 112308 287605
rect 112788 2619 112968 287605
rect 113448 2619 113628 287605
rect 114108 2619 127008 287605
rect 127488 2619 127668 287605
rect 128148 2619 128328 287605
rect 128808 2619 128988 287605
rect 129468 2619 142368 287605
rect 142848 2619 143028 287605
rect 143508 2619 143688 287605
rect 144168 2619 144348 287605
rect 144828 2619 157728 287605
rect 158208 2619 158388 287605
rect 158868 2619 159048 287605
rect 159528 2619 159708 287605
rect 160188 2619 173088 287605
rect 173568 2619 173748 287605
rect 174228 2619 174408 287605
rect 174888 2619 175068 287605
rect 175548 2619 188448 287605
rect 188928 2619 189108 287605
rect 189588 2619 189768 287605
rect 190248 2619 190428 287605
rect 190908 2619 203808 287605
rect 204288 2619 204468 287605
rect 204948 2619 205128 287605
rect 205608 2619 205788 287605
rect 206268 2619 219168 287605
rect 219648 2619 219828 287605
rect 220308 2619 220488 287605
rect 220968 2619 221148 287605
rect 221628 2619 234528 287605
rect 235008 2619 235188 287605
rect 235668 2619 235848 287605
rect 236328 2619 236508 287605
rect 236988 2619 249888 287605
rect 250368 2619 250548 287605
rect 251028 2619 251208 287605
rect 251688 2619 251868 287605
rect 252348 2619 265248 287605
rect 265728 2619 265908 287605
rect 266388 2619 266568 287605
rect 267048 2619 267228 287605
rect 267708 2619 280608 287605
rect 281088 2619 281268 287605
rect 281748 2619 281928 287605
rect 282408 2619 282588 287605
rect 283068 2619 283669 287605
<< labels >>
rlabel metal2 s 1214 289200 1270 290000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 76194 289200 76250 290000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 83646 289200 83702 290000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 91190 289200 91246 290000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 98642 289200 98698 290000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 106186 289200 106242 290000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 113638 289200 113694 290000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 121182 289200 121238 290000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 128634 289200 128690 290000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 136178 289200 136234 290000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 143630 289200 143686 290000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 8666 289200 8722 290000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 151174 289200 151230 290000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 158626 289200 158682 290000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 166170 289200 166226 290000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 173622 289200 173678 290000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 181166 289200 181222 290000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 188618 289200 188674 290000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 196162 289200 196218 290000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 203614 289200 203670 290000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 211158 289200 211214 290000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 218702 289200 218758 290000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 16210 289200 16266 290000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 226154 289200 226210 290000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 233698 289200 233754 290000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 241150 289200 241206 290000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 248694 289200 248750 290000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 256146 289200 256202 290000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 263690 289200 263746 290000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 271142 289200 271198 290000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 278686 289200 278742 290000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 23662 289200 23718 290000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 31206 289200 31262 290000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 38658 289200 38714 290000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 46202 289200 46258 290000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 53654 289200 53710 290000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 61198 289200 61254 290000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 68650 289200 68706 290000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3698 289200 3754 290000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 78678 289200 78734 290000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 86130 289200 86186 290000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 93674 289200 93730 290000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 101126 289200 101182 290000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 108670 289200 108726 290000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 116122 289200 116178 290000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 123666 289200 123722 290000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 131118 289200 131174 290000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 138662 289200 138718 290000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 146206 289200 146262 290000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 11150 289200 11206 290000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 153658 289200 153714 290000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 161202 289200 161258 290000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 168654 289200 168710 290000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 176198 289200 176254 290000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 183650 289200 183706 290000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 191194 289200 191250 290000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 198646 289200 198702 290000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 206190 289200 206246 290000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 213642 289200 213698 290000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 221186 289200 221242 290000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 18694 289200 18750 290000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 228638 289200 228694 290000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 236182 289200 236238 290000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 243634 289200 243690 290000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 251178 289200 251234 290000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 258630 289200 258686 290000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 266174 289200 266230 290000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 273626 289200 273682 290000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 281170 289200 281226 290000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 26146 289200 26202 290000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 33690 289200 33746 290000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 41142 289200 41198 290000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 48686 289200 48742 290000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 56138 289200 56194 290000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 63682 289200 63738 290000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 71134 289200 71190 290000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 6182 289200 6238 290000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 81162 289200 81218 290000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 88706 289200 88762 290000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 96158 289200 96214 290000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 103702 289200 103758 290000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 111154 289200 111210 290000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 118698 289200 118754 290000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 126150 289200 126206 290000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 133694 289200 133750 290000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 141146 289200 141202 290000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 148690 289200 148746 290000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 13634 289200 13690 290000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 156142 289200 156198 290000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 163686 289200 163742 290000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 171138 289200 171194 290000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 178682 289200 178738 290000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 186134 289200 186190 290000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 193678 289200 193734 290000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 201130 289200 201186 290000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 208674 289200 208730 290000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 216126 289200 216182 290000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 223670 289200 223726 290000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 21178 289200 21234 290000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 231122 289200 231178 290000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 238666 289200 238722 290000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 246118 289200 246174 290000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 253662 289200 253718 290000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 261114 289200 261170 290000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 268658 289200 268714 290000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 276110 289200 276166 290000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 283654 289200 283710 290000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 28630 289200 28686 290000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 36174 289200 36230 290000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 43626 289200 43682 290000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 51170 289200 51226 290000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 58622 289200 58678 290000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 66166 289200 66222 290000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 73710 289200 73766 290000 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 0 217472 800 217592 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 286138 289200 286194 290000 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 288622 289200 288678 290000 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 240506 0 240562 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 242254 0 242310 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 244094 0 244150 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 245842 0 245898 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 247590 0 247646 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 249430 0 249486 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 251178 0 251234 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 252926 0 252982 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 254766 0 254822 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 256514 0 256570 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 258262 0 258318 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 260010 0 260066 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 261850 0 261906 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 263598 0 263654 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 265346 0 265402 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 267186 0 267242 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 268934 0 268990 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 270682 0 270738 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 272522 0 272578 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 274270 0 274326 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 276018 0 276074 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 277766 0 277822 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 279606 0 279662 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 281354 0 281410 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 283102 0 283158 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 284942 0 284998 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 286690 0 286746 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 288438 0 288494 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 114466 0 114522 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 123298 0 123354 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 128634 0 128690 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 135810 0 135866 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 139306 0 139362 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 142894 0 142950 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 144642 0 144698 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 148230 0 148286 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 155314 0 155370 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 157062 0 157118 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 158810 0 158866 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 160650 0 160706 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 162398 0 162454 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 164146 0 164202 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 165986 0 166042 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 167734 0 167790 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 169482 0 169538 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 173070 0 173126 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 174818 0 174874 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 176566 0 176622 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 178406 0 178462 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 180154 0 180210 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 181902 0 181958 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 183742 0 183798 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 185490 0 185546 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 187238 0 187294 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 189078 0 189134 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 190826 0 190882 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 192574 0 192630 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 194322 0 194378 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 196162 0 196218 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 197910 0 197966 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 199658 0 199714 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 201498 0 201554 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 203246 0 203302 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 204994 0 205050 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 206742 0 206798 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 208582 0 208638 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 210330 0 210386 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 212078 0 212134 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 213918 0 213974 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 215666 0 215722 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 217414 0 217470 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 219254 0 219310 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 221002 0 221058 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 222750 0 222806 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 224498 0 224554 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 226338 0 226394 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 228086 0 228142 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 229834 0 229890 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 231674 0 231730 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 233422 0 233478 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 235170 0 235226 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 237010 0 237066 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 238758 0 238814 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 241150 0 241206 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 242898 0 242954 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 244646 0 244702 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 246394 0 246450 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 248234 0 248290 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 249982 0 250038 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 251730 0 251786 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 253570 0 253626 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 255318 0 255374 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 257066 0 257122 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 81346 0 81402 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 258906 0 258962 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 260654 0 260710 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 262402 0 262458 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 264150 0 264206 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 265990 0 266046 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 267738 0 267794 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 269486 0 269542 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 271326 0 271382 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 273074 0 273130 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 274822 0 274878 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 276662 0 276718 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 278410 0 278466 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 280158 0 280214 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 281906 0 281962 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 283746 0 283802 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 285494 0 285550 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 287242 0 287298 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 289082 0 289138 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 84842 0 84898 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 86682 0 86738 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 88430 0 88486 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 92018 0 92074 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 93766 0 93822 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 95514 0 95570 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 99102 0 99158 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 102598 0 102654 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 106186 0 106242 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 109774 0 109830 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 111522 0 111578 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 113270 0 113326 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 115018 0 115074 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 116858 0 116914 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 118606 0 118662 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 120354 0 120410 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 122194 0 122250 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 123942 0 123998 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 125690 0 125746 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 129278 0 129334 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 131026 0 131082 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 132774 0 132830 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 136362 0 136418 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 138110 0 138166 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 139950 0 140006 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 141698 0 141754 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 143446 0 143502 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 145286 0 145342 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 147034 0 147090 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 148782 0 148838 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 150530 0 150586 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 70674 0 70730 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 152370 0 152426 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 154118 0 154174 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 157706 0 157762 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 159454 0 159510 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 161202 0 161258 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 162950 0 163006 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 164790 0 164846 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 166538 0 166594 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 168286 0 168342 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 72422 0 72478 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 170126 0 170182 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 171874 0 171930 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 173622 0 173678 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 175462 0 175518 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 177210 0 177266 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 178958 0 179014 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 180706 0 180762 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 182546 0 182602 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 184294 0 184350 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 186042 0 186098 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 187882 0 187938 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 189630 0 189686 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 191378 0 191434 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 193218 0 193274 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 194966 0 195022 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 196714 0 196770 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 198462 0 198518 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 200302 0 200358 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 202050 0 202106 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 203798 0 203854 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 205638 0 205694 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 207386 0 207442 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 209134 0 209190 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 210974 0 211030 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 212722 0 212778 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 214470 0 214526 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 216218 0 216274 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 218058 0 218114 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 219806 0 219862 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 221554 0 221610 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 223394 0 223450 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 225142 0 225198 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 226890 0 226946 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 228730 0 228786 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 230478 0 230534 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 232226 0 232282 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 233974 0 234030 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 235814 0 235870 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 237562 0 237618 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 239310 0 239366 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 79506 0 79562 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 241702 0 241758 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 243450 0 243506 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 245290 0 245346 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 247038 0 247094 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 248786 0 248842 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 250626 0 250682 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 252374 0 252430 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 254122 0 254178 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 255870 0 255926 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 257710 0 257766 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 259458 0 259514 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 261206 0 261262 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 263046 0 263102 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 264794 0 264850 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 266542 0 266598 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 268290 0 268346 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 270130 0 270186 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 271878 0 271934 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 273626 0 273682 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 275466 0 275522 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 277214 0 277270 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 278962 0 279018 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 280802 0 280858 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 282550 0 282606 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 284298 0 284354 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 286046 0 286102 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 287886 0 287942 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 289634 0 289690 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 120998 0 121054 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 122746 0 122802 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 129830 0 129886 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 131670 0 131726 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 136914 0 136970 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 144090 0 144146 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 147586 0 147642 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 149426 0 149482 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 154670 0 154726 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 156510 0 156566 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 158258 0 158314 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 160006 0 160062 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 165342 0 165398 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 167182 0 167238 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 168930 0 168986 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 170678 0 170734 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 172426 0 172482 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 176014 0 176070 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 179602 0 179658 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 181350 0 181406 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 183098 0 183154 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 184846 0 184902 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 186686 0 186742 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 188434 0 188490 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 190182 0 190238 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 192022 0 192078 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 193770 0 193826 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 195518 0 195574 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 197358 0 197414 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 199106 0 199162 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 200854 0 200910 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 202602 0 202658 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 204442 0 204498 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 206190 0 206246 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 207938 0 207994 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 209778 0 209834 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 211526 0 211582 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 213274 0 213330 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 215114 0 215170 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 216862 0 216918 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 218610 0 218666 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 220358 0 220414 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 222198 0 222254 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 223946 0 224002 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 225694 0 225750 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 227534 0 227590 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 229282 0 229338 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 231030 0 231086 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 232870 0 232926 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 234618 0 234674 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 236366 0 236422 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 238114 0 238170 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 239954 0 240010 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal3 s 0 72496 800 72616 6 user_clk
port 502 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 503 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 504 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_ack_o
port 505 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 wbs_adr_i[0]
port 506 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_adr_i[10]
port 507 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_adr_i[11]
port 508 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wbs_adr_i[12]
port 509 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_adr_i[13]
port 510 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_adr_i[14]
port 511 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_adr_i[15]
port 512 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wbs_adr_i[16]
port 513 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_adr_i[17]
port 514 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 wbs_adr_i[18]
port 515 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 wbs_adr_i[19]
port 516 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_adr_i[1]
port 517 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 wbs_adr_i[20]
port 518 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 wbs_adr_i[21]
port 519 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 wbs_adr_i[22]
port 520 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 wbs_adr_i[23]
port 521 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 wbs_adr_i[24]
port 522 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 wbs_adr_i[25]
port 523 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 wbs_adr_i[26]
port 524 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 wbs_adr_i[27]
port 525 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 wbs_adr_i[28]
port 526 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 wbs_adr_i[29]
port 527 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_adr_i[2]
port 528 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 wbs_adr_i[30]
port 529 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 wbs_adr_i[31]
port 530 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_adr_i[3]
port 531 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_adr_i[4]
port 532 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_adr_i[5]
port 533 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_adr_i[6]
port 534 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[7]
port 535 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[8]
port 536 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_adr_i[9]
port 537 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_cyc_i
port 538 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_i[0]
port 539 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_dat_i[10]
port 540 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_dat_i[11]
port 541 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_i[12]
port 542 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 wbs_dat_i[13]
port 543 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_i[14]
port 544 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wbs_dat_i[15]
port 545 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wbs_dat_i[16]
port 546 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_i[17]
port 547 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 wbs_dat_i[18]
port 548 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_dat_i[19]
port 549 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_i[1]
port 550 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 wbs_dat_i[20]
port 551 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 wbs_dat_i[21]
port 552 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 wbs_dat_i[22]
port 553 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 wbs_dat_i[23]
port 554 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 wbs_dat_i[24]
port 555 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 wbs_dat_i[25]
port 556 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 wbs_dat_i[26]
port 557 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 wbs_dat_i[27]
port 558 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 wbs_dat_i[28]
port 559 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 wbs_dat_i[29]
port 560 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_dat_i[2]
port 561 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 wbs_dat_i[30]
port 562 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 wbs_dat_i[31]
port 563 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_i[3]
port 564 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[4]
port 565 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[5]
port 566 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_i[6]
port 567 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_dat_i[7]
port 568 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_i[8]
port 569 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_dat_i[9]
port 570 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_o[0]
port 571 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_o[10]
port 572 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_o[11]
port 573 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_o[12]
port 574 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_o[13]
port 575 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_o[14]
port 576 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_o[15]
port 577 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 wbs_dat_o[16]
port 578 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 wbs_dat_o[17]
port 579 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 wbs_dat_o[18]
port 580 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 wbs_dat_o[19]
port 581 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[1]
port 582 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 wbs_dat_o[20]
port 583 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 wbs_dat_o[21]
port 584 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 wbs_dat_o[22]
port 585 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 wbs_dat_o[23]
port 586 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 wbs_dat_o[24]
port 587 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 wbs_dat_o[25]
port 588 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 wbs_dat_o[26]
port 589 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 wbs_dat_o[27]
port 590 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 wbs_dat_o[28]
port 591 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 wbs_dat_o[29]
port 592 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_o[2]
port 593 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 wbs_dat_o[30]
port 594 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 wbs_dat_o[31]
port 595 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_o[3]
port 596 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_o[4]
port 597 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_o[5]
port 598 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 wbs_dat_o[6]
port 599 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_o[7]
port 600 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_o[8]
port 601 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_o[9]
port 602 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wbs_sel_i[0]
port 603 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_sel_i[1]
port 604 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_sel_i[2]
port 605 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_sel_i[3]
port 606 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_stb_i
port 607 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_we_i
port 608 nsew signal input
rlabel metal4 s 280688 2128 281008 287824 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 287824 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 287824 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 287824 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 287824 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 287824 6 vccd1
port 614 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 287824 6 vccd1
port 615 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 287824 6 vccd1
port 616 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 287824 6 vccd1
port 617 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 287824 6 vccd1
port 618 nsew power bidirectional
rlabel metal4 s 265328 2128 265648 287824 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 287824 6 vssd1
port 620 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 287824 6 vssd1
port 621 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 287824 6 vssd1
port 622 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 287824 6 vssd1
port 623 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 287824 6 vssd1
port 624 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 287824 6 vssd1
port 625 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 287824 6 vssd1
port 626 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 287824 6 vssd1
port 627 nsew ground bidirectional
rlabel metal4 s 281348 2176 281668 287776 6 vccd2
port 628 nsew power bidirectional
rlabel metal4 s 250628 2176 250948 287776 6 vccd2
port 629 nsew power bidirectional
rlabel metal4 s 219908 2176 220228 287776 6 vccd2
port 630 nsew power bidirectional
rlabel metal4 s 189188 2176 189508 287776 6 vccd2
port 631 nsew power bidirectional
rlabel metal4 s 158468 2176 158788 287776 6 vccd2
port 632 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 287776 6 vccd2
port 633 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 287776 6 vccd2
port 634 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 287776 6 vccd2
port 635 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 287776 6 vccd2
port 636 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 287776 6 vccd2
port 637 nsew power bidirectional
rlabel metal4 s 265988 2176 266308 287776 6 vssd2
port 638 nsew ground bidirectional
rlabel metal4 s 235268 2176 235588 287776 6 vssd2
port 639 nsew ground bidirectional
rlabel metal4 s 204548 2176 204868 287776 6 vssd2
port 640 nsew ground bidirectional
rlabel metal4 s 173828 2176 174148 287776 6 vssd2
port 641 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 287776 6 vssd2
port 642 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 287776 6 vssd2
port 643 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 287776 6 vssd2
port 644 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 287776 6 vssd2
port 645 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 287776 6 vssd2
port 646 nsew ground bidirectional
rlabel metal4 s 282008 2176 282328 287776 6 vdda1
port 647 nsew power bidirectional
rlabel metal4 s 251288 2176 251608 287776 6 vdda1
port 648 nsew power bidirectional
rlabel metal4 s 220568 2176 220888 287776 6 vdda1
port 649 nsew power bidirectional
rlabel metal4 s 189848 2176 190168 287776 6 vdda1
port 650 nsew power bidirectional
rlabel metal4 s 159128 2176 159448 287776 6 vdda1
port 651 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 287776 6 vdda1
port 652 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 287776 6 vdda1
port 653 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 287776 6 vdda1
port 654 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 287776 6 vdda1
port 655 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 287776 6 vdda1
port 656 nsew power bidirectional
rlabel metal4 s 266648 2176 266968 287776 6 vssa1
port 657 nsew ground bidirectional
rlabel metal4 s 235928 2176 236248 287776 6 vssa1
port 658 nsew ground bidirectional
rlabel metal4 s 205208 2176 205528 287776 6 vssa1
port 659 nsew ground bidirectional
rlabel metal4 s 174488 2176 174808 287776 6 vssa1
port 660 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 287776 6 vssa1
port 661 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 287776 6 vssa1
port 662 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 287776 6 vssa1
port 663 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 287776 6 vssa1
port 664 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 287776 6 vssa1
port 665 nsew ground bidirectional
rlabel metal4 s 282668 2176 282988 287776 6 vdda2
port 666 nsew power bidirectional
rlabel metal4 s 251948 2176 252268 287776 6 vdda2
port 667 nsew power bidirectional
rlabel metal4 s 221228 2176 221548 287776 6 vdda2
port 668 nsew power bidirectional
rlabel metal4 s 190508 2176 190828 287776 6 vdda2
port 669 nsew power bidirectional
rlabel metal4 s 159788 2176 160108 287776 6 vdda2
port 670 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 287776 6 vdda2
port 671 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 287776 6 vdda2
port 672 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 287776 6 vdda2
port 673 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 287776 6 vdda2
port 674 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 287776 6 vdda2
port 675 nsew power bidirectional
rlabel metal4 s 267308 2176 267628 287776 6 vssa2
port 676 nsew ground bidirectional
rlabel metal4 s 236588 2176 236908 287776 6 vssa2
port 677 nsew ground bidirectional
rlabel metal4 s 205868 2176 206188 287776 6 vssa2
port 678 nsew ground bidirectional
rlabel metal4 s 175148 2176 175468 287776 6 vssa2
port 679 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 287776 6 vssa2
port 680 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 287776 6 vssa2
port 681 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 287776 6 vssa2
port 682 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 287776 6 vssa2
port 683 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 287776 6 vssa2
port 684 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 290000 290000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 262967018
string GDS_START 853434
<< end >>

