magic
tech sky130A
magscale 1 2
timestamp 1623069705
<< obsli1 >>
rect 1104 2159 198812 197489
<< obsm1 >>
rect 198 1368 199810 197520
<< metal2 >>
rect 846 199200 902 200000
rect 2502 199200 2558 200000
rect 4250 199200 4306 200000
rect 5998 199200 6054 200000
rect 7746 199200 7802 200000
rect 9494 199200 9550 200000
rect 11242 199200 11298 200000
rect 12990 199200 13046 200000
rect 14738 199200 14794 200000
rect 16486 199200 16542 200000
rect 18234 199200 18290 200000
rect 19890 199200 19946 200000
rect 21638 199200 21694 200000
rect 23386 199200 23442 200000
rect 25134 199200 25190 200000
rect 26882 199200 26938 200000
rect 28630 199200 28686 200000
rect 30378 199200 30434 200000
rect 32126 199200 32182 200000
rect 33874 199200 33930 200000
rect 35622 199200 35678 200000
rect 37278 199200 37334 200000
rect 39026 199200 39082 200000
rect 40774 199200 40830 200000
rect 42522 199200 42578 200000
rect 44270 199200 44326 200000
rect 46018 199200 46074 200000
rect 47766 199200 47822 200000
rect 49514 199200 49570 200000
rect 51262 199200 51318 200000
rect 53010 199200 53066 200000
rect 54758 199200 54814 200000
rect 56414 199200 56470 200000
rect 58162 199200 58218 200000
rect 59910 199200 59966 200000
rect 61658 199200 61714 200000
rect 63406 199200 63462 200000
rect 65154 199200 65210 200000
rect 66902 199200 66958 200000
rect 68650 199200 68706 200000
rect 70398 199200 70454 200000
rect 72146 199200 72202 200000
rect 73802 199200 73858 200000
rect 75550 199200 75606 200000
rect 77298 199200 77354 200000
rect 79046 199200 79102 200000
rect 80794 199200 80850 200000
rect 82542 199200 82598 200000
rect 84290 199200 84346 200000
rect 86038 199200 86094 200000
rect 87786 199200 87842 200000
rect 89534 199200 89590 200000
rect 91282 199200 91338 200000
rect 92938 199200 92994 200000
rect 94686 199200 94742 200000
rect 96434 199200 96490 200000
rect 98182 199200 98238 200000
rect 99930 199200 99986 200000
rect 101678 199200 101734 200000
rect 103426 199200 103482 200000
rect 105174 199200 105230 200000
rect 106922 199200 106978 200000
rect 108670 199200 108726 200000
rect 110326 199200 110382 200000
rect 112074 199200 112130 200000
rect 113822 199200 113878 200000
rect 115570 199200 115626 200000
rect 117318 199200 117374 200000
rect 119066 199200 119122 200000
rect 120814 199200 120870 200000
rect 122562 199200 122618 200000
rect 124310 199200 124366 200000
rect 126058 199200 126114 200000
rect 127806 199200 127862 200000
rect 129462 199200 129518 200000
rect 131210 199200 131266 200000
rect 132958 199200 133014 200000
rect 134706 199200 134762 200000
rect 136454 199200 136510 200000
rect 138202 199200 138258 200000
rect 139950 199200 140006 200000
rect 141698 199200 141754 200000
rect 143446 199200 143502 200000
rect 145194 199200 145250 200000
rect 146850 199200 146906 200000
rect 148598 199200 148654 200000
rect 150346 199200 150402 200000
rect 152094 199200 152150 200000
rect 153842 199200 153898 200000
rect 155590 199200 155646 200000
rect 157338 199200 157394 200000
rect 159086 199200 159142 200000
rect 160834 199200 160890 200000
rect 162582 199200 162638 200000
rect 164330 199200 164386 200000
rect 165986 199200 166042 200000
rect 167734 199200 167790 200000
rect 169482 199200 169538 200000
rect 171230 199200 171286 200000
rect 172978 199200 173034 200000
rect 174726 199200 174782 200000
rect 176474 199200 176530 200000
rect 178222 199200 178278 200000
rect 179970 199200 180026 200000
rect 181718 199200 181774 200000
rect 183374 199200 183430 200000
rect 185122 199200 185178 200000
rect 186870 199200 186926 200000
rect 188618 199200 188674 200000
rect 190366 199200 190422 200000
rect 192114 199200 192170 200000
rect 193862 199200 193918 200000
rect 195610 199200 195666 200000
rect 197358 199200 197414 200000
rect 199106 199200 199162 200000
rect 202 0 258 800
rect 570 0 626 800
rect 938 0 994 800
rect 1398 0 1454 800
rect 1766 0 1822 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 3054 0 3110 800
rect 3422 0 3478 800
rect 3790 0 3846 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 5078 0 5134 800
rect 5446 0 5502 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7102 0 7158 800
rect 7470 0 7526 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8758 0 8814 800
rect 9126 0 9182 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10782 0 10838 800
rect 11150 0 11206 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12438 0 12494 800
rect 12806 0 12862 800
rect 13174 0 13230 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18142 0 18198 800
rect 18510 0 18566 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20166 0 20222 800
rect 20534 0 20590 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21822 0 21878 800
rect 22190 0 22246 800
rect 22650 0 22706 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23846 0 23902 800
rect 24214 0 24270 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25502 0 25558 800
rect 25870 0 25926 800
rect 26238 0 26294 800
rect 26698 0 26754 800
rect 27066 0 27122 800
rect 27526 0 27582 800
rect 27894 0 27950 800
rect 28354 0 28410 800
rect 28722 0 28778 800
rect 29182 0 29238 800
rect 29550 0 29606 800
rect 29918 0 29974 800
rect 30378 0 30434 800
rect 30746 0 30802 800
rect 31206 0 31262 800
rect 31574 0 31630 800
rect 32034 0 32090 800
rect 32402 0 32458 800
rect 32770 0 32826 800
rect 33230 0 33286 800
rect 33598 0 33654 800
rect 34058 0 34114 800
rect 34426 0 34482 800
rect 34886 0 34942 800
rect 35254 0 35310 800
rect 35622 0 35678 800
rect 36082 0 36138 800
rect 36450 0 36506 800
rect 36910 0 36966 800
rect 37278 0 37334 800
rect 37738 0 37794 800
rect 38106 0 38162 800
rect 38566 0 38622 800
rect 38934 0 38990 800
rect 39302 0 39358 800
rect 39762 0 39818 800
rect 40130 0 40186 800
rect 40590 0 40646 800
rect 40958 0 41014 800
rect 41418 0 41474 800
rect 41786 0 41842 800
rect 42154 0 42210 800
rect 42614 0 42670 800
rect 42982 0 43038 800
rect 43442 0 43498 800
rect 43810 0 43866 800
rect 44270 0 44326 800
rect 44638 0 44694 800
rect 45098 0 45154 800
rect 45466 0 45522 800
rect 45834 0 45890 800
rect 46294 0 46350 800
rect 46662 0 46718 800
rect 47122 0 47178 800
rect 47490 0 47546 800
rect 47950 0 48006 800
rect 48318 0 48374 800
rect 48686 0 48742 800
rect 49146 0 49202 800
rect 49514 0 49570 800
rect 49974 0 50030 800
rect 50342 0 50398 800
rect 50802 0 50858 800
rect 51170 0 51226 800
rect 51630 0 51686 800
rect 51998 0 52054 800
rect 52366 0 52422 800
rect 52826 0 52882 800
rect 53194 0 53250 800
rect 53654 0 53710 800
rect 54022 0 54078 800
rect 54482 0 54538 800
rect 54850 0 54906 800
rect 55218 0 55274 800
rect 55678 0 55734 800
rect 56046 0 56102 800
rect 56506 0 56562 800
rect 56874 0 56930 800
rect 57334 0 57390 800
rect 57702 0 57758 800
rect 58162 0 58218 800
rect 58530 0 58586 800
rect 58898 0 58954 800
rect 59358 0 59414 800
rect 59726 0 59782 800
rect 60186 0 60242 800
rect 60554 0 60610 800
rect 61014 0 61070 800
rect 61382 0 61438 800
rect 61750 0 61806 800
rect 62210 0 62266 800
rect 62578 0 62634 800
rect 63038 0 63094 800
rect 63406 0 63462 800
rect 63866 0 63922 800
rect 64234 0 64290 800
rect 64694 0 64750 800
rect 65062 0 65118 800
rect 65430 0 65486 800
rect 65890 0 65946 800
rect 66258 0 66314 800
rect 66718 0 66774 800
rect 67086 0 67142 800
rect 67546 0 67602 800
rect 67914 0 67970 800
rect 68282 0 68338 800
rect 68742 0 68798 800
rect 69110 0 69166 800
rect 69570 0 69626 800
rect 69938 0 69994 800
rect 70398 0 70454 800
rect 70766 0 70822 800
rect 71134 0 71190 800
rect 71594 0 71650 800
rect 71962 0 72018 800
rect 72422 0 72478 800
rect 72790 0 72846 800
rect 73250 0 73306 800
rect 73618 0 73674 800
rect 74078 0 74134 800
rect 74446 0 74502 800
rect 74814 0 74870 800
rect 75274 0 75330 800
rect 75642 0 75698 800
rect 76102 0 76158 800
rect 76470 0 76526 800
rect 76930 0 76986 800
rect 77298 0 77354 800
rect 77666 0 77722 800
rect 78126 0 78182 800
rect 78494 0 78550 800
rect 78954 0 79010 800
rect 79322 0 79378 800
rect 79782 0 79838 800
rect 80150 0 80206 800
rect 80610 0 80666 800
rect 80978 0 81034 800
rect 81346 0 81402 800
rect 81806 0 81862 800
rect 82174 0 82230 800
rect 82634 0 82690 800
rect 83002 0 83058 800
rect 83462 0 83518 800
rect 83830 0 83886 800
rect 84198 0 84254 800
rect 84658 0 84714 800
rect 85026 0 85082 800
rect 85486 0 85542 800
rect 85854 0 85910 800
rect 86314 0 86370 800
rect 86682 0 86738 800
rect 87142 0 87198 800
rect 87510 0 87566 800
rect 87878 0 87934 800
rect 88338 0 88394 800
rect 88706 0 88762 800
rect 89166 0 89222 800
rect 89534 0 89590 800
rect 89994 0 90050 800
rect 90362 0 90418 800
rect 90730 0 90786 800
rect 91190 0 91246 800
rect 91558 0 91614 800
rect 92018 0 92074 800
rect 92386 0 92442 800
rect 92846 0 92902 800
rect 93214 0 93270 800
rect 93674 0 93730 800
rect 94042 0 94098 800
rect 94410 0 94466 800
rect 94870 0 94926 800
rect 95238 0 95294 800
rect 95698 0 95754 800
rect 96066 0 96122 800
rect 96526 0 96582 800
rect 96894 0 96950 800
rect 97262 0 97318 800
rect 97722 0 97778 800
rect 98090 0 98146 800
rect 98550 0 98606 800
rect 98918 0 98974 800
rect 99378 0 99434 800
rect 99746 0 99802 800
rect 100206 0 100262 800
rect 100574 0 100630 800
rect 100942 0 100998 800
rect 101402 0 101458 800
rect 101770 0 101826 800
rect 102230 0 102286 800
rect 102598 0 102654 800
rect 103058 0 103114 800
rect 103426 0 103482 800
rect 103794 0 103850 800
rect 104254 0 104310 800
rect 104622 0 104678 800
rect 105082 0 105138 800
rect 105450 0 105506 800
rect 105910 0 105966 800
rect 106278 0 106334 800
rect 106646 0 106702 800
rect 107106 0 107162 800
rect 107474 0 107530 800
rect 107934 0 107990 800
rect 108302 0 108358 800
rect 108762 0 108818 800
rect 109130 0 109186 800
rect 109590 0 109646 800
rect 109958 0 110014 800
rect 110326 0 110382 800
rect 110786 0 110842 800
rect 111154 0 111210 800
rect 111614 0 111670 800
rect 111982 0 112038 800
rect 112442 0 112498 800
rect 112810 0 112866 800
rect 113178 0 113234 800
rect 113638 0 113694 800
rect 114006 0 114062 800
rect 114466 0 114522 800
rect 114834 0 114890 800
rect 115294 0 115350 800
rect 115662 0 115718 800
rect 116122 0 116178 800
rect 116490 0 116546 800
rect 116858 0 116914 800
rect 117318 0 117374 800
rect 117686 0 117742 800
rect 118146 0 118202 800
rect 118514 0 118570 800
rect 118974 0 119030 800
rect 119342 0 119398 800
rect 119710 0 119766 800
rect 120170 0 120226 800
rect 120538 0 120594 800
rect 120998 0 121054 800
rect 121366 0 121422 800
rect 121826 0 121882 800
rect 122194 0 122250 800
rect 122654 0 122710 800
rect 123022 0 123078 800
rect 123390 0 123446 800
rect 123850 0 123906 800
rect 124218 0 124274 800
rect 124678 0 124734 800
rect 125046 0 125102 800
rect 125506 0 125562 800
rect 125874 0 125930 800
rect 126242 0 126298 800
rect 126702 0 126758 800
rect 127070 0 127126 800
rect 127530 0 127586 800
rect 127898 0 127954 800
rect 128358 0 128414 800
rect 128726 0 128782 800
rect 129186 0 129242 800
rect 129554 0 129610 800
rect 129922 0 129978 800
rect 130382 0 130438 800
rect 130750 0 130806 800
rect 131210 0 131266 800
rect 131578 0 131634 800
rect 132038 0 132094 800
rect 132406 0 132462 800
rect 132774 0 132830 800
rect 133234 0 133290 800
rect 133602 0 133658 800
rect 134062 0 134118 800
rect 134430 0 134486 800
rect 134890 0 134946 800
rect 135258 0 135314 800
rect 135626 0 135682 800
rect 136086 0 136142 800
rect 136454 0 136510 800
rect 136914 0 136970 800
rect 137282 0 137338 800
rect 137742 0 137798 800
rect 138110 0 138166 800
rect 138570 0 138626 800
rect 138938 0 138994 800
rect 139306 0 139362 800
rect 139766 0 139822 800
rect 140134 0 140190 800
rect 140594 0 140650 800
rect 140962 0 141018 800
rect 141422 0 141478 800
rect 141790 0 141846 800
rect 142158 0 142214 800
rect 142618 0 142674 800
rect 142986 0 143042 800
rect 143446 0 143502 800
rect 143814 0 143870 800
rect 144274 0 144330 800
rect 144642 0 144698 800
rect 145102 0 145158 800
rect 145470 0 145526 800
rect 145838 0 145894 800
rect 146298 0 146354 800
rect 146666 0 146722 800
rect 147126 0 147182 800
rect 147494 0 147550 800
rect 147954 0 148010 800
rect 148322 0 148378 800
rect 148690 0 148746 800
rect 149150 0 149206 800
rect 149518 0 149574 800
rect 149978 0 150034 800
rect 150346 0 150402 800
rect 150806 0 150862 800
rect 151174 0 151230 800
rect 151634 0 151690 800
rect 152002 0 152058 800
rect 152370 0 152426 800
rect 152830 0 152886 800
rect 153198 0 153254 800
rect 153658 0 153714 800
rect 154026 0 154082 800
rect 154486 0 154542 800
rect 154854 0 154910 800
rect 155222 0 155278 800
rect 155682 0 155738 800
rect 156050 0 156106 800
rect 156510 0 156566 800
rect 156878 0 156934 800
rect 157338 0 157394 800
rect 157706 0 157762 800
rect 158166 0 158222 800
rect 158534 0 158590 800
rect 158902 0 158958 800
rect 159362 0 159418 800
rect 159730 0 159786 800
rect 160190 0 160246 800
rect 160558 0 160614 800
rect 161018 0 161074 800
rect 161386 0 161442 800
rect 161754 0 161810 800
rect 162214 0 162270 800
rect 162582 0 162638 800
rect 163042 0 163098 800
rect 163410 0 163466 800
rect 163870 0 163926 800
rect 164238 0 164294 800
rect 164698 0 164754 800
rect 165066 0 165122 800
rect 165434 0 165490 800
rect 165894 0 165950 800
rect 166262 0 166318 800
rect 166722 0 166778 800
rect 167090 0 167146 800
rect 167550 0 167606 800
rect 167918 0 167974 800
rect 168286 0 168342 800
rect 168746 0 168802 800
rect 169114 0 169170 800
rect 169574 0 169630 800
rect 169942 0 169998 800
rect 170402 0 170458 800
rect 170770 0 170826 800
rect 171138 0 171194 800
rect 171598 0 171654 800
rect 171966 0 172022 800
rect 172426 0 172482 800
rect 172794 0 172850 800
rect 173254 0 173310 800
rect 173622 0 173678 800
rect 174082 0 174138 800
rect 174450 0 174506 800
rect 174818 0 174874 800
rect 175278 0 175334 800
rect 175646 0 175702 800
rect 176106 0 176162 800
rect 176474 0 176530 800
rect 176934 0 176990 800
rect 177302 0 177358 800
rect 177670 0 177726 800
rect 178130 0 178186 800
rect 178498 0 178554 800
rect 178958 0 179014 800
rect 179326 0 179382 800
rect 179786 0 179842 800
rect 180154 0 180210 800
rect 180614 0 180670 800
rect 180982 0 181038 800
rect 181350 0 181406 800
rect 181810 0 181866 800
rect 182178 0 182234 800
rect 182638 0 182694 800
rect 183006 0 183062 800
rect 183466 0 183522 800
rect 183834 0 183890 800
rect 184202 0 184258 800
rect 184662 0 184718 800
rect 185030 0 185086 800
rect 185490 0 185546 800
rect 185858 0 185914 800
rect 186318 0 186374 800
rect 186686 0 186742 800
rect 187146 0 187202 800
rect 187514 0 187570 800
rect 187882 0 187938 800
rect 188342 0 188398 800
rect 188710 0 188766 800
rect 189170 0 189226 800
rect 189538 0 189594 800
rect 189998 0 190054 800
rect 190366 0 190422 800
rect 190734 0 190790 800
rect 191194 0 191250 800
rect 191562 0 191618 800
rect 192022 0 192078 800
rect 192390 0 192446 800
rect 192850 0 192906 800
rect 193218 0 193274 800
rect 193678 0 193734 800
rect 194046 0 194102 800
rect 194414 0 194470 800
rect 194874 0 194930 800
rect 195242 0 195298 800
rect 195702 0 195758 800
rect 196070 0 196126 800
rect 196530 0 196586 800
rect 196898 0 196954 800
rect 197266 0 197322 800
rect 197726 0 197782 800
rect 198094 0 198150 800
rect 198554 0 198610 800
rect 198922 0 198978 800
rect 199382 0 199438 800
rect 199750 0 199806 800
<< obsm2 >>
rect 204 199144 790 199200
rect 958 199144 2446 199200
rect 2614 199144 4194 199200
rect 4362 199144 5942 199200
rect 6110 199144 7690 199200
rect 7858 199144 9438 199200
rect 9606 199144 11186 199200
rect 11354 199144 12934 199200
rect 13102 199144 14682 199200
rect 14850 199144 16430 199200
rect 16598 199144 18178 199200
rect 18346 199144 19834 199200
rect 20002 199144 21582 199200
rect 21750 199144 23330 199200
rect 23498 199144 25078 199200
rect 25246 199144 26826 199200
rect 26994 199144 28574 199200
rect 28742 199144 30322 199200
rect 30490 199144 32070 199200
rect 32238 199144 33818 199200
rect 33986 199144 35566 199200
rect 35734 199144 37222 199200
rect 37390 199144 38970 199200
rect 39138 199144 40718 199200
rect 40886 199144 42466 199200
rect 42634 199144 44214 199200
rect 44382 199144 45962 199200
rect 46130 199144 47710 199200
rect 47878 199144 49458 199200
rect 49626 199144 51206 199200
rect 51374 199144 52954 199200
rect 53122 199144 54702 199200
rect 54870 199144 56358 199200
rect 56526 199144 58106 199200
rect 58274 199144 59854 199200
rect 60022 199144 61602 199200
rect 61770 199144 63350 199200
rect 63518 199144 65098 199200
rect 65266 199144 66846 199200
rect 67014 199144 68594 199200
rect 68762 199144 70342 199200
rect 70510 199144 72090 199200
rect 72258 199144 73746 199200
rect 73914 199144 75494 199200
rect 75662 199144 77242 199200
rect 77410 199144 78990 199200
rect 79158 199144 80738 199200
rect 80906 199144 82486 199200
rect 82654 199144 84234 199200
rect 84402 199144 85982 199200
rect 86150 199144 87730 199200
rect 87898 199144 89478 199200
rect 89646 199144 91226 199200
rect 91394 199144 92882 199200
rect 93050 199144 94630 199200
rect 94798 199144 96378 199200
rect 96546 199144 98126 199200
rect 98294 199144 99874 199200
rect 100042 199144 101622 199200
rect 101790 199144 103370 199200
rect 103538 199144 105118 199200
rect 105286 199144 106866 199200
rect 107034 199144 108614 199200
rect 108782 199144 110270 199200
rect 110438 199144 112018 199200
rect 112186 199144 113766 199200
rect 113934 199144 115514 199200
rect 115682 199144 117262 199200
rect 117430 199144 119010 199200
rect 119178 199144 120758 199200
rect 120926 199144 122506 199200
rect 122674 199144 124254 199200
rect 124422 199144 126002 199200
rect 126170 199144 127750 199200
rect 127918 199144 129406 199200
rect 129574 199144 131154 199200
rect 131322 199144 132902 199200
rect 133070 199144 134650 199200
rect 134818 199144 136398 199200
rect 136566 199144 138146 199200
rect 138314 199144 139894 199200
rect 140062 199144 141642 199200
rect 141810 199144 143390 199200
rect 143558 199144 145138 199200
rect 145306 199144 146794 199200
rect 146962 199144 148542 199200
rect 148710 199144 150290 199200
rect 150458 199144 152038 199200
rect 152206 199144 153786 199200
rect 153954 199144 155534 199200
rect 155702 199144 157282 199200
rect 157450 199144 159030 199200
rect 159198 199144 160778 199200
rect 160946 199144 162526 199200
rect 162694 199144 164274 199200
rect 164442 199144 165930 199200
rect 166098 199144 167678 199200
rect 167846 199144 169426 199200
rect 169594 199144 171174 199200
rect 171342 199144 172922 199200
rect 173090 199144 174670 199200
rect 174838 199144 176418 199200
rect 176586 199144 178166 199200
rect 178334 199144 179914 199200
rect 180082 199144 181662 199200
rect 181830 199144 183318 199200
rect 183486 199144 185066 199200
rect 185234 199144 186814 199200
rect 186982 199144 188562 199200
rect 188730 199144 190310 199200
rect 190478 199144 192058 199200
rect 192226 199144 193806 199200
rect 193974 199144 195554 199200
rect 195722 199144 197302 199200
rect 197470 199144 199050 199200
rect 199218 199144 199804 199200
rect 204 856 199804 199144
rect 314 800 514 856
rect 682 800 882 856
rect 1050 800 1342 856
rect 1510 800 1710 856
rect 1878 800 2170 856
rect 2338 800 2538 856
rect 2706 800 2998 856
rect 3166 800 3366 856
rect 3534 800 3734 856
rect 3902 800 4194 856
rect 4362 800 4562 856
rect 4730 800 5022 856
rect 5190 800 5390 856
rect 5558 800 5850 856
rect 6018 800 6218 856
rect 6386 800 6586 856
rect 6754 800 7046 856
rect 7214 800 7414 856
rect 7582 800 7874 856
rect 8042 800 8242 856
rect 8410 800 8702 856
rect 8870 800 9070 856
rect 9238 800 9530 856
rect 9698 800 9898 856
rect 10066 800 10266 856
rect 10434 800 10726 856
rect 10894 800 11094 856
rect 11262 800 11554 856
rect 11722 800 11922 856
rect 12090 800 12382 856
rect 12550 800 12750 856
rect 12918 800 13118 856
rect 13286 800 13578 856
rect 13746 800 13946 856
rect 14114 800 14406 856
rect 14574 800 14774 856
rect 14942 800 15234 856
rect 15402 800 15602 856
rect 15770 800 16062 856
rect 16230 800 16430 856
rect 16598 800 16798 856
rect 16966 800 17258 856
rect 17426 800 17626 856
rect 17794 800 18086 856
rect 18254 800 18454 856
rect 18622 800 18914 856
rect 19082 800 19282 856
rect 19450 800 19650 856
rect 19818 800 20110 856
rect 20278 800 20478 856
rect 20646 800 20938 856
rect 21106 800 21306 856
rect 21474 800 21766 856
rect 21934 800 22134 856
rect 22302 800 22594 856
rect 22762 800 22962 856
rect 23130 800 23330 856
rect 23498 800 23790 856
rect 23958 800 24158 856
rect 24326 800 24618 856
rect 24786 800 24986 856
rect 25154 800 25446 856
rect 25614 800 25814 856
rect 25982 800 26182 856
rect 26350 800 26642 856
rect 26810 800 27010 856
rect 27178 800 27470 856
rect 27638 800 27838 856
rect 28006 800 28298 856
rect 28466 800 28666 856
rect 28834 800 29126 856
rect 29294 800 29494 856
rect 29662 800 29862 856
rect 30030 800 30322 856
rect 30490 800 30690 856
rect 30858 800 31150 856
rect 31318 800 31518 856
rect 31686 800 31978 856
rect 32146 800 32346 856
rect 32514 800 32714 856
rect 32882 800 33174 856
rect 33342 800 33542 856
rect 33710 800 34002 856
rect 34170 800 34370 856
rect 34538 800 34830 856
rect 34998 800 35198 856
rect 35366 800 35566 856
rect 35734 800 36026 856
rect 36194 800 36394 856
rect 36562 800 36854 856
rect 37022 800 37222 856
rect 37390 800 37682 856
rect 37850 800 38050 856
rect 38218 800 38510 856
rect 38678 800 38878 856
rect 39046 800 39246 856
rect 39414 800 39706 856
rect 39874 800 40074 856
rect 40242 800 40534 856
rect 40702 800 40902 856
rect 41070 800 41362 856
rect 41530 800 41730 856
rect 41898 800 42098 856
rect 42266 800 42558 856
rect 42726 800 42926 856
rect 43094 800 43386 856
rect 43554 800 43754 856
rect 43922 800 44214 856
rect 44382 800 44582 856
rect 44750 800 45042 856
rect 45210 800 45410 856
rect 45578 800 45778 856
rect 45946 800 46238 856
rect 46406 800 46606 856
rect 46774 800 47066 856
rect 47234 800 47434 856
rect 47602 800 47894 856
rect 48062 800 48262 856
rect 48430 800 48630 856
rect 48798 800 49090 856
rect 49258 800 49458 856
rect 49626 800 49918 856
rect 50086 800 50286 856
rect 50454 800 50746 856
rect 50914 800 51114 856
rect 51282 800 51574 856
rect 51742 800 51942 856
rect 52110 800 52310 856
rect 52478 800 52770 856
rect 52938 800 53138 856
rect 53306 800 53598 856
rect 53766 800 53966 856
rect 54134 800 54426 856
rect 54594 800 54794 856
rect 54962 800 55162 856
rect 55330 800 55622 856
rect 55790 800 55990 856
rect 56158 800 56450 856
rect 56618 800 56818 856
rect 56986 800 57278 856
rect 57446 800 57646 856
rect 57814 800 58106 856
rect 58274 800 58474 856
rect 58642 800 58842 856
rect 59010 800 59302 856
rect 59470 800 59670 856
rect 59838 800 60130 856
rect 60298 800 60498 856
rect 60666 800 60958 856
rect 61126 800 61326 856
rect 61494 800 61694 856
rect 61862 800 62154 856
rect 62322 800 62522 856
rect 62690 800 62982 856
rect 63150 800 63350 856
rect 63518 800 63810 856
rect 63978 800 64178 856
rect 64346 800 64638 856
rect 64806 800 65006 856
rect 65174 800 65374 856
rect 65542 800 65834 856
rect 66002 800 66202 856
rect 66370 800 66662 856
rect 66830 800 67030 856
rect 67198 800 67490 856
rect 67658 800 67858 856
rect 68026 800 68226 856
rect 68394 800 68686 856
rect 68854 800 69054 856
rect 69222 800 69514 856
rect 69682 800 69882 856
rect 70050 800 70342 856
rect 70510 800 70710 856
rect 70878 800 71078 856
rect 71246 800 71538 856
rect 71706 800 71906 856
rect 72074 800 72366 856
rect 72534 800 72734 856
rect 72902 800 73194 856
rect 73362 800 73562 856
rect 73730 800 74022 856
rect 74190 800 74390 856
rect 74558 800 74758 856
rect 74926 800 75218 856
rect 75386 800 75586 856
rect 75754 800 76046 856
rect 76214 800 76414 856
rect 76582 800 76874 856
rect 77042 800 77242 856
rect 77410 800 77610 856
rect 77778 800 78070 856
rect 78238 800 78438 856
rect 78606 800 78898 856
rect 79066 800 79266 856
rect 79434 800 79726 856
rect 79894 800 80094 856
rect 80262 800 80554 856
rect 80722 800 80922 856
rect 81090 800 81290 856
rect 81458 800 81750 856
rect 81918 800 82118 856
rect 82286 800 82578 856
rect 82746 800 82946 856
rect 83114 800 83406 856
rect 83574 800 83774 856
rect 83942 800 84142 856
rect 84310 800 84602 856
rect 84770 800 84970 856
rect 85138 800 85430 856
rect 85598 800 85798 856
rect 85966 800 86258 856
rect 86426 800 86626 856
rect 86794 800 87086 856
rect 87254 800 87454 856
rect 87622 800 87822 856
rect 87990 800 88282 856
rect 88450 800 88650 856
rect 88818 800 89110 856
rect 89278 800 89478 856
rect 89646 800 89938 856
rect 90106 800 90306 856
rect 90474 800 90674 856
rect 90842 800 91134 856
rect 91302 800 91502 856
rect 91670 800 91962 856
rect 92130 800 92330 856
rect 92498 800 92790 856
rect 92958 800 93158 856
rect 93326 800 93618 856
rect 93786 800 93986 856
rect 94154 800 94354 856
rect 94522 800 94814 856
rect 94982 800 95182 856
rect 95350 800 95642 856
rect 95810 800 96010 856
rect 96178 800 96470 856
rect 96638 800 96838 856
rect 97006 800 97206 856
rect 97374 800 97666 856
rect 97834 800 98034 856
rect 98202 800 98494 856
rect 98662 800 98862 856
rect 99030 800 99322 856
rect 99490 800 99690 856
rect 99858 800 100150 856
rect 100318 800 100518 856
rect 100686 800 100886 856
rect 101054 800 101346 856
rect 101514 800 101714 856
rect 101882 800 102174 856
rect 102342 800 102542 856
rect 102710 800 103002 856
rect 103170 800 103370 856
rect 103538 800 103738 856
rect 103906 800 104198 856
rect 104366 800 104566 856
rect 104734 800 105026 856
rect 105194 800 105394 856
rect 105562 800 105854 856
rect 106022 800 106222 856
rect 106390 800 106590 856
rect 106758 800 107050 856
rect 107218 800 107418 856
rect 107586 800 107878 856
rect 108046 800 108246 856
rect 108414 800 108706 856
rect 108874 800 109074 856
rect 109242 800 109534 856
rect 109702 800 109902 856
rect 110070 800 110270 856
rect 110438 800 110730 856
rect 110898 800 111098 856
rect 111266 800 111558 856
rect 111726 800 111926 856
rect 112094 800 112386 856
rect 112554 800 112754 856
rect 112922 800 113122 856
rect 113290 800 113582 856
rect 113750 800 113950 856
rect 114118 800 114410 856
rect 114578 800 114778 856
rect 114946 800 115238 856
rect 115406 800 115606 856
rect 115774 800 116066 856
rect 116234 800 116434 856
rect 116602 800 116802 856
rect 116970 800 117262 856
rect 117430 800 117630 856
rect 117798 800 118090 856
rect 118258 800 118458 856
rect 118626 800 118918 856
rect 119086 800 119286 856
rect 119454 800 119654 856
rect 119822 800 120114 856
rect 120282 800 120482 856
rect 120650 800 120942 856
rect 121110 800 121310 856
rect 121478 800 121770 856
rect 121938 800 122138 856
rect 122306 800 122598 856
rect 122766 800 122966 856
rect 123134 800 123334 856
rect 123502 800 123794 856
rect 123962 800 124162 856
rect 124330 800 124622 856
rect 124790 800 124990 856
rect 125158 800 125450 856
rect 125618 800 125818 856
rect 125986 800 126186 856
rect 126354 800 126646 856
rect 126814 800 127014 856
rect 127182 800 127474 856
rect 127642 800 127842 856
rect 128010 800 128302 856
rect 128470 800 128670 856
rect 128838 800 129130 856
rect 129298 800 129498 856
rect 129666 800 129866 856
rect 130034 800 130326 856
rect 130494 800 130694 856
rect 130862 800 131154 856
rect 131322 800 131522 856
rect 131690 800 131982 856
rect 132150 800 132350 856
rect 132518 800 132718 856
rect 132886 800 133178 856
rect 133346 800 133546 856
rect 133714 800 134006 856
rect 134174 800 134374 856
rect 134542 800 134834 856
rect 135002 800 135202 856
rect 135370 800 135570 856
rect 135738 800 136030 856
rect 136198 800 136398 856
rect 136566 800 136858 856
rect 137026 800 137226 856
rect 137394 800 137686 856
rect 137854 800 138054 856
rect 138222 800 138514 856
rect 138682 800 138882 856
rect 139050 800 139250 856
rect 139418 800 139710 856
rect 139878 800 140078 856
rect 140246 800 140538 856
rect 140706 800 140906 856
rect 141074 800 141366 856
rect 141534 800 141734 856
rect 141902 800 142102 856
rect 142270 800 142562 856
rect 142730 800 142930 856
rect 143098 800 143390 856
rect 143558 800 143758 856
rect 143926 800 144218 856
rect 144386 800 144586 856
rect 144754 800 145046 856
rect 145214 800 145414 856
rect 145582 800 145782 856
rect 145950 800 146242 856
rect 146410 800 146610 856
rect 146778 800 147070 856
rect 147238 800 147438 856
rect 147606 800 147898 856
rect 148066 800 148266 856
rect 148434 800 148634 856
rect 148802 800 149094 856
rect 149262 800 149462 856
rect 149630 800 149922 856
rect 150090 800 150290 856
rect 150458 800 150750 856
rect 150918 800 151118 856
rect 151286 800 151578 856
rect 151746 800 151946 856
rect 152114 800 152314 856
rect 152482 800 152774 856
rect 152942 800 153142 856
rect 153310 800 153602 856
rect 153770 800 153970 856
rect 154138 800 154430 856
rect 154598 800 154798 856
rect 154966 800 155166 856
rect 155334 800 155626 856
rect 155794 800 155994 856
rect 156162 800 156454 856
rect 156622 800 156822 856
rect 156990 800 157282 856
rect 157450 800 157650 856
rect 157818 800 158110 856
rect 158278 800 158478 856
rect 158646 800 158846 856
rect 159014 800 159306 856
rect 159474 800 159674 856
rect 159842 800 160134 856
rect 160302 800 160502 856
rect 160670 800 160962 856
rect 161130 800 161330 856
rect 161498 800 161698 856
rect 161866 800 162158 856
rect 162326 800 162526 856
rect 162694 800 162986 856
rect 163154 800 163354 856
rect 163522 800 163814 856
rect 163982 800 164182 856
rect 164350 800 164642 856
rect 164810 800 165010 856
rect 165178 800 165378 856
rect 165546 800 165838 856
rect 166006 800 166206 856
rect 166374 800 166666 856
rect 166834 800 167034 856
rect 167202 800 167494 856
rect 167662 800 167862 856
rect 168030 800 168230 856
rect 168398 800 168690 856
rect 168858 800 169058 856
rect 169226 800 169518 856
rect 169686 800 169886 856
rect 170054 800 170346 856
rect 170514 800 170714 856
rect 170882 800 171082 856
rect 171250 800 171542 856
rect 171710 800 171910 856
rect 172078 800 172370 856
rect 172538 800 172738 856
rect 172906 800 173198 856
rect 173366 800 173566 856
rect 173734 800 174026 856
rect 174194 800 174394 856
rect 174562 800 174762 856
rect 174930 800 175222 856
rect 175390 800 175590 856
rect 175758 800 176050 856
rect 176218 800 176418 856
rect 176586 800 176878 856
rect 177046 800 177246 856
rect 177414 800 177614 856
rect 177782 800 178074 856
rect 178242 800 178442 856
rect 178610 800 178902 856
rect 179070 800 179270 856
rect 179438 800 179730 856
rect 179898 800 180098 856
rect 180266 800 180558 856
rect 180726 800 180926 856
rect 181094 800 181294 856
rect 181462 800 181754 856
rect 181922 800 182122 856
rect 182290 800 182582 856
rect 182750 800 182950 856
rect 183118 800 183410 856
rect 183578 800 183778 856
rect 183946 800 184146 856
rect 184314 800 184606 856
rect 184774 800 184974 856
rect 185142 800 185434 856
rect 185602 800 185802 856
rect 185970 800 186262 856
rect 186430 800 186630 856
rect 186798 800 187090 856
rect 187258 800 187458 856
rect 187626 800 187826 856
rect 187994 800 188286 856
rect 188454 800 188654 856
rect 188822 800 189114 856
rect 189282 800 189482 856
rect 189650 800 189942 856
rect 190110 800 190310 856
rect 190478 800 190678 856
rect 190846 800 191138 856
rect 191306 800 191506 856
rect 191674 800 191966 856
rect 192134 800 192334 856
rect 192502 800 192794 856
rect 192962 800 193162 856
rect 193330 800 193622 856
rect 193790 800 193990 856
rect 194158 800 194358 856
rect 194526 800 194818 856
rect 194986 800 195186 856
rect 195354 800 195646 856
rect 195814 800 196014 856
rect 196182 800 196474 856
rect 196642 800 196842 856
rect 197010 800 197210 856
rect 197378 800 197670 856
rect 197838 800 198038 856
rect 198206 800 198498 856
rect 198666 800 198866 856
rect 199034 800 199326 856
rect 199494 800 199694 856
<< metal3 >>
rect 0 99968 800 100088
rect 199200 99968 200000 100088
<< obsm3 >>
rect 800 100168 199200 197505
rect 880 99888 199120 100168
rect 800 2143 199200 99888
<< metal4 >>
rect 4208 2128 4528 197520
rect 4868 2176 5188 197472
rect 5528 2176 5848 197472
rect 6188 2176 6508 197472
rect 19568 2128 19888 197520
rect 20228 2176 20548 197472
rect 20888 2176 21208 197472
rect 21548 2176 21868 197472
rect 34928 2128 35248 197520
rect 35588 2176 35908 197472
rect 36248 2176 36568 197472
rect 36908 2176 37228 197472
rect 50288 2128 50608 197520
rect 50948 2176 51268 197472
rect 51608 2176 51928 197472
rect 52268 2176 52588 197472
rect 65648 2128 65968 197520
rect 66308 2176 66628 197472
rect 66968 2176 67288 197472
rect 67628 2176 67948 197472
rect 81008 2128 81328 197520
rect 81668 2176 81988 197472
rect 82328 2176 82648 197472
rect 82988 2176 83308 197472
rect 96368 2128 96688 197520
rect 97028 2176 97348 197472
rect 97688 2176 98008 197472
rect 98348 2176 98668 197472
rect 111728 2128 112048 197520
rect 112388 2176 112708 197472
rect 113048 2176 113368 197472
rect 113708 2176 114028 197472
rect 127088 2128 127408 197520
rect 127748 2176 128068 197472
rect 128408 2176 128728 197472
rect 129068 2176 129388 197472
rect 142448 2128 142768 197520
rect 143108 2176 143428 197472
rect 143768 2176 144088 197472
rect 144428 2176 144748 197472
rect 157808 2128 158128 197520
rect 158468 2176 158788 197472
rect 159128 2176 159448 197472
rect 159788 2176 160108 197472
rect 173168 2128 173488 197520
rect 173828 2176 174148 197472
rect 174488 2176 174808 197472
rect 175148 2176 175468 197472
rect 188528 2128 188848 197520
rect 189188 2176 189508 197472
rect 189848 2176 190168 197472
rect 190508 2176 190828 197472
<< obsm4 >>
rect 84331 41243 96288 121413
rect 96768 41243 96948 121413
rect 97428 41243 97608 121413
rect 98088 41243 98268 121413
rect 98748 41243 111648 121413
rect 112128 41243 112308 121413
rect 112788 41243 112968 121413
rect 113448 41243 113628 121413
rect 114108 41243 127008 121413
rect 127488 41243 127668 121413
rect 128148 41243 128328 121413
rect 128808 41243 128988 121413
rect 129468 41243 142368 121413
rect 142848 41243 143028 121413
rect 143508 41243 143688 121413
rect 144168 41243 144348 121413
rect 144828 41243 157728 121413
rect 158208 41243 158388 121413
rect 158868 41243 159048 121413
rect 159528 41243 159708 121413
rect 160188 41243 164069 121413
<< labels >>
rlabel metal2 s 846 199200 902 200000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 53010 199200 53066 200000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 58162 199200 58218 200000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 63406 199200 63462 200000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 68650 199200 68706 200000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 73802 199200 73858 200000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 79046 199200 79102 200000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 84290 199200 84346 200000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 89534 199200 89590 200000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 94686 199200 94742 200000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 99930 199200 99986 200000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5998 199200 6054 200000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 105174 199200 105230 200000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 110326 199200 110382 200000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 115570 199200 115626 200000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 120814 199200 120870 200000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 126058 199200 126114 200000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 131210 199200 131266 200000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 136454 199200 136510 200000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 141698 199200 141754 200000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 146850 199200 146906 200000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 152094 199200 152150 200000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 11242 199200 11298 200000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 157338 199200 157394 200000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 162582 199200 162638 200000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 167734 199200 167790 200000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 172978 199200 173034 200000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 178222 199200 178278 200000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 183374 199200 183430 200000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 188618 199200 188674 200000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 193862 199200 193918 200000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 16486 199200 16542 200000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 21638 199200 21694 200000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 26882 199200 26938 200000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 32126 199200 32182 200000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 37278 199200 37334 200000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 42522 199200 42578 200000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 47766 199200 47822 200000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2502 199200 2558 200000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 54758 199200 54814 200000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 59910 199200 59966 200000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 65154 199200 65210 200000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 70398 199200 70454 200000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 75550 199200 75606 200000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 80794 199200 80850 200000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 86038 199200 86094 200000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 91282 199200 91338 200000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 96434 199200 96490 200000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 101678 199200 101734 200000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7746 199200 7802 200000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 106922 199200 106978 200000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 112074 199200 112130 200000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 117318 199200 117374 200000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 122562 199200 122618 200000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 127806 199200 127862 200000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 132958 199200 133014 200000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 138202 199200 138258 200000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 143446 199200 143502 200000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 148598 199200 148654 200000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 153842 199200 153898 200000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 12990 199200 13046 200000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 159086 199200 159142 200000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 164330 199200 164386 200000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 169482 199200 169538 200000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 174726 199200 174782 200000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 179970 199200 180026 200000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 185122 199200 185178 200000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 190366 199200 190422 200000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 195610 199200 195666 200000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 18234 199200 18290 200000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 23386 199200 23442 200000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 28630 199200 28686 200000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 33874 199200 33930 200000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 39026 199200 39082 200000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 44270 199200 44326 200000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 49514 199200 49570 200000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4250 199200 4306 200000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 56414 199200 56470 200000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 61658 199200 61714 200000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 66902 199200 66958 200000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 72146 199200 72202 200000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 77298 199200 77354 200000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 82542 199200 82598 200000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 87786 199200 87842 200000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 92938 199200 92994 200000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 98182 199200 98238 200000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 103426 199200 103482 200000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 9494 199200 9550 200000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 108670 199200 108726 200000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 113822 199200 113878 200000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 119066 199200 119122 200000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 124310 199200 124366 200000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 129462 199200 129518 200000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 134706 199200 134762 200000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 139950 199200 140006 200000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 145194 199200 145250 200000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 150346 199200 150402 200000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 155590 199200 155646 200000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 14738 199200 14794 200000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 160834 199200 160890 200000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 165986 199200 166042 200000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 171230 199200 171286 200000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 176474 199200 176530 200000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 181718 199200 181774 200000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 186870 199200 186926 200000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 192114 199200 192170 200000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 197358 199200 197414 200000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 19890 199200 19946 200000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 25134 199200 25190 200000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 30378 199200 30434 200000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 35622 199200 35678 200000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 40774 199200 40830 200000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 46018 199200 46074 200000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 51262 199200 51318 200000 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 199200 99968 200000 100088 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 199106 199200 199162 200000 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 165894 0 165950 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 167090 0 167146 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 168286 0 168342 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 169574 0 169630 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 170770 0 170826 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 171966 0 172022 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 173254 0 173310 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 174450 0 174506 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 175646 0 175702 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 176934 0 176990 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 178130 0 178186 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 179326 0 179382 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 180614 0 180670 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 181810 0 181866 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 183006 0 183062 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 184202 0 184258 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 185490 0 185546 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 186686 0 186742 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 187882 0 187938 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 189170 0 189226 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 190366 0 190422 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 191562 0 191618 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 192850 0 192906 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 194046 0 194102 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 195242 0 195298 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 196530 0 196586 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 197726 0 197782 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 198922 0 198978 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 114466 0 114522 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 121826 0 121882 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 124218 0 124274 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 126702 0 126758 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 132774 0 132830 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 137742 0 137798 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 140134 0 140190 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 141422 0 141478 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 152370 0 152426 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 156050 0 156106 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 158534 0 158590 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 162214 0 162270 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 163410 0 163466 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 166262 0 166318 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 167550 0 167606 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 168746 0 168802 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 169942 0 169998 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 171138 0 171194 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 172426 0 172482 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 173622 0 173678 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 174818 0 174874 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 176106 0 176162 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 177302 0 177358 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 178498 0 178554 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 179786 0 179842 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 180982 0 181038 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 182178 0 182234 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 183466 0 183522 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 184662 0 184718 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 185858 0 185914 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 187146 0 187202 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 188342 0 188398 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 189538 0 189594 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 190734 0 190790 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 192022 0 192078 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 193218 0 193274 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 194414 0 194470 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 195702 0 195758 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 196898 0 196954 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 198094 0 198150 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 199382 0 199438 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 61014 0 61070 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 71962 0 72018 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 73250 0 73306 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 76930 0 76986 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 79322 0 79378 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 83002 0 83058 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 84198 0 84254 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 85486 0 85542 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 86682 0 86738 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 90362 0 90418 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 47490 0 47546 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 92846 0 92902 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 95238 0 95294 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 96526 0 96582 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 97722 0 97778 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 101402 0 101458 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 102598 0 102654 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 103794 0 103850 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 105082 0 105138 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 107474 0 107530 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 108762 0 108818 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 109958 0 110014 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 111154 0 111210 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 112442 0 112498 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 114834 0 114890 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 116122 0 116178 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 117318 0 117374 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 119710 0 119766 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 120998 0 121054 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 122194 0 122250 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 123390 0 123446 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 124678 0 124734 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 125874 0 125930 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 127070 0 127126 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 128358 0 128414 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 51170 0 51226 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 129554 0 129610 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 133234 0 133290 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 134430 0 134486 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 135626 0 135682 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 136914 0 136970 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 138110 0 138166 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 139306 0 139362 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 140594 0 140650 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 52366 0 52422 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 141790 0 141846 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 142986 0 143042 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 144274 0 144330 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 145470 0 145526 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 146666 0 146722 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 147954 0 148010 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 149150 0 149206 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 150346 0 150402 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 151634 0 151690 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 152830 0 152886 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 154026 0 154082 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 155222 0 155278 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 156510 0 156566 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 157706 0 157762 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 158902 0 158958 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 160190 0 160246 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 161386 0 161442 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 162582 0 162638 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 165066 0 165122 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 54850 0 54906 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 166722 0 166778 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 167918 0 167974 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 170402 0 170458 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 171598 0 171654 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 172794 0 172850 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 174082 0 174138 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 175278 0 175334 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 177670 0 177726 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 178958 0 179014 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 180154 0 180210 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 181350 0 181406 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 183834 0 183890 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 185030 0 185086 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 186318 0 186374 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 187514 0 187570 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 188710 0 188766 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 191194 0 191250 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 192390 0 192446 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 193678 0 193734 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 194874 0 194930 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 196070 0 196126 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 197266 0 197322 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 198554 0 198610 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 199750 0 199806 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 106646 0 106702 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 125046 0 125102 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 132406 0 132462 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 136086 0 136142 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 138570 0 138626 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 139766 0 139822 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 140962 0 141018 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 143446 0 143502 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 144642 0 144698 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 147126 0 147182 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 150806 0 150862 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 154486 0 154542 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 155682 0 155738 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 158166 0 158222 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 159362 0 159418 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 160558 0 160614 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 161754 0 161810 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 163042 0 163098 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 164238 0 164294 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 165434 0 165490 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 570 0 626 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_ack_o
port 504 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_dat_o[0]
port 570 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_o[10]
port 571 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_o[11]
port 572 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_o[12]
port 573 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_o[13]
port 574 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_o[14]
port 575 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[15]
port 576 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_o[16]
port 577 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 wbs_dat_o[17]
port 578 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 wbs_dat_o[18]
port 579 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_o[19]
port 580 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_o[1]
port 581 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 wbs_dat_o[20]
port 582 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_o[21]
port 583 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[22]
port 584 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_o[23]
port 585 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 wbs_dat_o[24]
port 586 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 wbs_dat_o[25]
port 587 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_o[26]
port 588 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 wbs_dat_o[27]
port 589 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 wbs_dat_o[28]
port 590 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 wbs_dat_o[29]
port 591 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 wbs_dat_o[2]
port 592 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 wbs_dat_o[30]
port 593 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 wbs_dat_o[31]
port 594 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_o[3]
port 595 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[4]
port 596 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_o[5]
port 597 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_o[6]
port 598 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_o[7]
port 599 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[8]
port 600 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_o[9]
port 601 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 188528 2128 188848 197520 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 197520 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 197520 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 197520 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 197520 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 614 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 197520 6 vssd1
port 615 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 197520 6 vssd1
port 616 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 197520 6 vssd1
port 617 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 197520 6 vssd1
port 618 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 197520 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 620 nsew ground bidirectional
rlabel metal4 s 189188 2176 189508 197472 6 vccd2
port 621 nsew power bidirectional
rlabel metal4 s 158468 2176 158788 197472 6 vccd2
port 622 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 197472 6 vccd2
port 623 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 197472 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 197472 6 vccd2
port 625 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 197472 6 vccd2
port 626 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 197472 6 vccd2
port 627 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 197472 6 vssd2
port 628 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 197472 6 vssd2
port 629 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 197472 6 vssd2
port 630 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 197472 6 vssd2
port 631 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 197472 6 vssd2
port 632 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 197472 6 vssd2
port 633 nsew ground bidirectional
rlabel metal4 s 189848 2176 190168 197472 6 vdda1
port 634 nsew power bidirectional
rlabel metal4 s 159128 2176 159448 197472 6 vdda1
port 635 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 197472 6 vdda1
port 636 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 197472 6 vdda1
port 637 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 197472 6 vdda1
port 638 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 197472 6 vdda1
port 639 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 197472 6 vdda1
port 640 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 197472 6 vssa1
port 641 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 197472 6 vssa1
port 642 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 197472 6 vssa1
port 643 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 197472 6 vssa1
port 644 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 197472 6 vssa1
port 645 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 197472 6 vssa1
port 646 nsew ground bidirectional
rlabel metal4 s 190508 2176 190828 197472 6 vdda2
port 647 nsew power bidirectional
rlabel metal4 s 159788 2176 160108 197472 6 vdda2
port 648 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 197472 6 vdda2
port 649 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 197472 6 vdda2
port 650 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 197472 6 vdda2
port 651 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 197472 6 vdda2
port 652 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 197472 6 vdda2
port 653 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 197472 6 vssa2
port 654 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 197472 6 vssa2
port 655 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 197472 6 vssa2
port 656 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 197472 6 vssa2
port 657 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 197472 6 vssa2
port 658 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 197472 6 vssa2
port 659 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 200000 200000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj.gds
string GDS_END 41003308
string GDS_START 795838
<< end >>

