`default_nettype none
//-----------------------------------------------------
// Project Name : a.out
// Function     : Main processor 
// Description  : This is the main processor
// Coder        : Jaquer AND VORIXO

//***Headers***

//***Module***
module state_counters #(
        parameter integer WORD_SIZE = 32,
        parameter integer VERIFICATION_PINS = 2,
        parameter integer WHISBONE_ADR = 32,
        parameter integer COUNTERSIZE = 32,
        parameter [31:0]  ADDRBASE     = 32'h3000_0000,
        parameter [31:0]  COUNTERDATA  = ADDRBASE + 4
    )
    (
        `ifdef USE_POWER_PINS
        inout vdda1,	// User area 1 3.3V supply
        inout vdda2,	// User area 2 3.3V supply
        inout vssa1,	// User area 1 analog ground
        inout vssa2,	// User area 2 analog ground
        inout vccd1,	// User area 1 1.8V supply
        inout vccd2,	// User area 2 1.8v supply
        inout vssd1,	// User area 1 digital ground
        inout vssd2,	// User area 2 digital ground
        `endif
        input  clk_i ,
        input  rst_i ,
        input  valid_i, 
        input  [3 : 0] wstrb_i,
        input  [WORD_SIZE -1 : 0] wdata_i,
        input  [WHISBONE_ADR - 1 : 0] whisbone_addr_i,
        input  [VERIFICATION_PINS - 1 : 0] operation_result_i ,
        input  valid_output_i,
        input  wbs_we_i,
        output  ready_o,
        output [WORD_SIZE - 1 : 0] rdata_o
    );

//***Internal logic generated by compiler***  


//***Dumped Internal logic***
    reg [COUNTERSIZE-1:0] ecc_corrected_errors;
    reg [COUNTERSIZE-1:0] ecc_uncorrected_errors;
    reg [COUNTERSIZE-1:0] total_reads;
    reg ready_o;
    reg [WORD_SIZE-1:0] rdata_o;


    always @(posedge clk_i) begin

        if(rst_i) begin
            total_reads <= {WORD_SIZE {1'b0}}; 
            ecc_uncorrected_errors <= {WORD_SIZE {1'b0}}; 
            ecc_corrected_errors <= {WORD_SIZE {1'b0}}; 
            ready_o <= 1'b0;
        end
        else begin
            if (valid_output_i == 1'b1) begin
                total_reads <= total_reads +1;
                if (operation_result_i[0] == 1'b1) begin
                    ecc_corrected_errors <= ecc_corrected_errors + 1;
                end
                if (operation_result_i[1] == 1'b1) begin
                    ecc_uncorrected_errors <= ecc_uncorrected_errors + 1;
                end
            end
            if (valid_i) begin
                case (whisbone_addr_i)
                COUNTERDATA : begin
                        ready_o <= 1'b1;
                        if (wbs_we_i) begin
                            if (wstrb_i[0]) total_reads[7:0]   <= wdata_i[7:0];
                            if (wstrb_i[1]) total_reads[15:8]  <= wdata_i[15:8];
                            if (wstrb_i[2]) total_reads[23:16] <= wdata_i[23:16];
                            if (wstrb_i[3]) total_reads[31:24] <= wdata_i[31:24];
                        end
                        else begin
                            rdata_o = total_reads;
                        end
                    end
                COUNTERDATA + 4: begin
                        ready_o <= 1'b1;
                        rdata_o = ecc_corrected_errors;
                        if (wbs_we_i) begin
                            if (wstrb_i[0]) ecc_corrected_errors[7:0]   <= wdata_i[7:0];
                            if (wstrb_i[1]) ecc_corrected_errors[15:8]  <= wdata_i[15:8];
                            if (wstrb_i[2]) ecc_corrected_errors[23:16] <= wdata_i[23:16];
                            if (wstrb_i[3]) ecc_corrected_errors[31:24] <= wdata_i[31:24];
                        end
                        else begin
                            rdata_o = ecc_corrected_errors;
                        end
                    end
                COUNTERDATA + 8: begin
                        ready_o <= 1'b1;
                        if (wbs_we_i) begin
                            if (wstrb_i[0]) ecc_uncorrected_errors[7:0]   <= wdata_i[7:0];
                            if (wstrb_i[1]) ecc_uncorrected_errors[15:8]  <= wdata_i[15:8];
                            if (wstrb_i[2]) ecc_uncorrected_errors[23:16] <= wdata_i[23:16];
                            if (wstrb_i[3]) ecc_uncorrected_errors[31:24] <= wdata_i[31:24];
                        end
                        else begin
                            rdata_o = ecc_uncorrected_errors;
                        end
                    end
                ADDRBASE: begin
                        ready_o <= 1'b1;
                    end
                default: ready_o <= 1'b0;
                
                endcase
                
            end
        end
    end

    
//***Handcrafted Internal logic*** 
//TODO
endmodule
