magic
tech sky130A
magscale 1 2
timestamp 1625592194
<< obsli1 >>
rect 1104 2159 297039 295409
<< obsm1 >>
rect 290 1164 297698 295440
<< metal2 >>
rect 1306 297200 1362 298000
rect 3882 297200 3938 298000
rect 6458 297200 6514 298000
rect 9126 297200 9182 298000
rect 11702 297200 11758 298000
rect 14370 297200 14426 298000
rect 16946 297200 17002 298000
rect 19522 297200 19578 298000
rect 22190 297200 22246 298000
rect 24766 297200 24822 298000
rect 27434 297200 27490 298000
rect 30010 297200 30066 298000
rect 32586 297200 32642 298000
rect 35254 297200 35310 298000
rect 37830 297200 37886 298000
rect 40498 297200 40554 298000
rect 43074 297200 43130 298000
rect 45742 297200 45798 298000
rect 48318 297200 48374 298000
rect 50894 297200 50950 298000
rect 53562 297200 53618 298000
rect 56138 297200 56194 298000
rect 58806 297200 58862 298000
rect 61382 297200 61438 298000
rect 63958 297200 64014 298000
rect 66626 297200 66682 298000
rect 69202 297200 69258 298000
rect 71870 297200 71926 298000
rect 74446 297200 74502 298000
rect 77022 297200 77078 298000
rect 79690 297200 79746 298000
rect 82266 297200 82322 298000
rect 84934 297200 84990 298000
rect 87510 297200 87566 298000
rect 90178 297200 90234 298000
rect 92754 297200 92810 298000
rect 95330 297200 95386 298000
rect 97998 297200 98054 298000
rect 100574 297200 100630 298000
rect 103242 297200 103298 298000
rect 105818 297200 105874 298000
rect 108394 297200 108450 298000
rect 111062 297200 111118 298000
rect 113638 297200 113694 298000
rect 116306 297200 116362 298000
rect 118882 297200 118938 298000
rect 121458 297200 121514 298000
rect 124126 297200 124182 298000
rect 126702 297200 126758 298000
rect 129370 297200 129426 298000
rect 131946 297200 132002 298000
rect 134614 297200 134670 298000
rect 137190 297200 137246 298000
rect 139766 297200 139822 298000
rect 142434 297200 142490 298000
rect 145010 297200 145066 298000
rect 147678 297200 147734 298000
rect 150254 297200 150310 298000
rect 152830 297200 152886 298000
rect 155498 297200 155554 298000
rect 158074 297200 158130 298000
rect 160742 297200 160798 298000
rect 163318 297200 163374 298000
rect 165894 297200 165950 298000
rect 168562 297200 168618 298000
rect 171138 297200 171194 298000
rect 173806 297200 173862 298000
rect 176382 297200 176438 298000
rect 179050 297200 179106 298000
rect 181626 297200 181682 298000
rect 184202 297200 184258 298000
rect 186870 297200 186926 298000
rect 189446 297200 189502 298000
rect 192114 297200 192170 298000
rect 194690 297200 194746 298000
rect 197266 297200 197322 298000
rect 199934 297200 199990 298000
rect 202510 297200 202566 298000
rect 205178 297200 205234 298000
rect 207754 297200 207810 298000
rect 210330 297200 210386 298000
rect 212998 297200 213054 298000
rect 215574 297200 215630 298000
rect 218242 297200 218298 298000
rect 220818 297200 220874 298000
rect 223486 297200 223542 298000
rect 226062 297200 226118 298000
rect 228638 297200 228694 298000
rect 231306 297200 231362 298000
rect 233882 297200 233938 298000
rect 236550 297200 236606 298000
rect 239126 297200 239182 298000
rect 241702 297200 241758 298000
rect 244370 297200 244426 298000
rect 246946 297200 247002 298000
rect 249614 297200 249670 298000
rect 252190 297200 252246 298000
rect 254766 297200 254822 298000
rect 257434 297200 257490 298000
rect 260010 297200 260066 298000
rect 262678 297200 262734 298000
rect 265254 297200 265310 298000
rect 267922 297200 267978 298000
rect 270498 297200 270554 298000
rect 273074 297200 273130 298000
rect 275742 297200 275798 298000
rect 278318 297200 278374 298000
rect 280986 297200 281042 298000
rect 283562 297200 283618 298000
rect 286138 297200 286194 298000
rect 288806 297200 288862 298000
rect 291382 297200 291438 298000
rect 294050 297200 294106 298000
rect 296626 297200 296682 298000
rect 294 0 350 800
rect 846 0 902 800
rect 1490 0 1546 800
rect 2042 0 2098 800
rect 2686 0 2742 800
rect 3330 0 3386 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5722 0 5778 800
rect 6366 0 6422 800
rect 6918 0 6974 800
rect 7562 0 7618 800
rect 8114 0 8170 800
rect 8758 0 8814 800
rect 9402 0 9458 800
rect 9954 0 10010 800
rect 10598 0 10654 800
rect 11150 0 11206 800
rect 11794 0 11850 800
rect 12438 0 12494 800
rect 12990 0 13046 800
rect 13634 0 13690 800
rect 14278 0 14334 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16026 0 16082 800
rect 16670 0 16726 800
rect 17314 0 17370 800
rect 17866 0 17922 800
rect 18510 0 18566 800
rect 19062 0 19118 800
rect 19706 0 19762 800
rect 20350 0 20406 800
rect 20902 0 20958 800
rect 21546 0 21602 800
rect 22098 0 22154 800
rect 22742 0 22798 800
rect 23386 0 23442 800
rect 23938 0 23994 800
rect 24582 0 24638 800
rect 25226 0 25282 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 26974 0 27030 800
rect 27618 0 27674 800
rect 28262 0 28318 800
rect 28814 0 28870 800
rect 29458 0 29514 800
rect 30010 0 30066 800
rect 30654 0 30710 800
rect 31298 0 31354 800
rect 31850 0 31906 800
rect 32494 0 32550 800
rect 33046 0 33102 800
rect 33690 0 33746 800
rect 34334 0 34390 800
rect 34886 0 34942 800
rect 35530 0 35586 800
rect 36174 0 36230 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 37922 0 37978 800
rect 38566 0 38622 800
rect 39210 0 39266 800
rect 39762 0 39818 800
rect 40406 0 40462 800
rect 40958 0 41014 800
rect 41602 0 41658 800
rect 42246 0 42302 800
rect 42798 0 42854 800
rect 43442 0 43498 800
rect 43994 0 44050 800
rect 44638 0 44694 800
rect 45282 0 45338 800
rect 45834 0 45890 800
rect 46478 0 46534 800
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 48870 0 48926 800
rect 49514 0 49570 800
rect 50158 0 50214 800
rect 50710 0 50766 800
rect 51354 0 51410 800
rect 51906 0 51962 800
rect 52550 0 52606 800
rect 53194 0 53250 800
rect 53746 0 53802 800
rect 54390 0 54446 800
rect 54942 0 54998 800
rect 55586 0 55642 800
rect 56230 0 56286 800
rect 56782 0 56838 800
rect 57426 0 57482 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 59818 0 59874 800
rect 60462 0 60518 800
rect 61106 0 61162 800
rect 61658 0 61714 800
rect 62302 0 62358 800
rect 62854 0 62910 800
rect 63498 0 63554 800
rect 64142 0 64198 800
rect 64694 0 64750 800
rect 65338 0 65394 800
rect 65890 0 65946 800
rect 66534 0 66590 800
rect 67178 0 67234 800
rect 67730 0 67786 800
rect 68374 0 68430 800
rect 68926 0 68982 800
rect 69570 0 69626 800
rect 70214 0 70270 800
rect 70766 0 70822 800
rect 71410 0 71466 800
rect 72054 0 72110 800
rect 72606 0 72662 800
rect 73250 0 73306 800
rect 73802 0 73858 800
rect 74446 0 74502 800
rect 75090 0 75146 800
rect 75642 0 75698 800
rect 76286 0 76342 800
rect 76838 0 76894 800
rect 77482 0 77538 800
rect 78126 0 78182 800
rect 78678 0 78734 800
rect 79322 0 79378 800
rect 79874 0 79930 800
rect 80518 0 80574 800
rect 81162 0 81218 800
rect 81714 0 81770 800
rect 82358 0 82414 800
rect 82910 0 82966 800
rect 83554 0 83610 800
rect 84198 0 84254 800
rect 84750 0 84806 800
rect 85394 0 85450 800
rect 86038 0 86094 800
rect 86590 0 86646 800
rect 87234 0 87290 800
rect 87786 0 87842 800
rect 88430 0 88486 800
rect 89074 0 89130 800
rect 89626 0 89682 800
rect 90270 0 90326 800
rect 90822 0 90878 800
rect 91466 0 91522 800
rect 92110 0 92166 800
rect 92662 0 92718 800
rect 93306 0 93362 800
rect 93858 0 93914 800
rect 94502 0 94558 800
rect 95146 0 95202 800
rect 95698 0 95754 800
rect 96342 0 96398 800
rect 96986 0 97042 800
rect 97538 0 97594 800
rect 98182 0 98238 800
rect 98734 0 98790 800
rect 99378 0 99434 800
rect 100022 0 100078 800
rect 100574 0 100630 800
rect 101218 0 101274 800
rect 101770 0 101826 800
rect 102414 0 102470 800
rect 103058 0 103114 800
rect 103610 0 103666 800
rect 104254 0 104310 800
rect 104806 0 104862 800
rect 105450 0 105506 800
rect 106094 0 106150 800
rect 106646 0 106702 800
rect 107290 0 107346 800
rect 107934 0 107990 800
rect 108486 0 108542 800
rect 109130 0 109186 800
rect 109682 0 109738 800
rect 110326 0 110382 800
rect 110970 0 111026 800
rect 111522 0 111578 800
rect 112166 0 112222 800
rect 112718 0 112774 800
rect 113362 0 113418 800
rect 114006 0 114062 800
rect 114558 0 114614 800
rect 115202 0 115258 800
rect 115754 0 115810 800
rect 116398 0 116454 800
rect 117042 0 117098 800
rect 117594 0 117650 800
rect 118238 0 118294 800
rect 118790 0 118846 800
rect 119434 0 119490 800
rect 120078 0 120134 800
rect 120630 0 120686 800
rect 121274 0 121330 800
rect 121918 0 121974 800
rect 122470 0 122526 800
rect 123114 0 123170 800
rect 123666 0 123722 800
rect 124310 0 124366 800
rect 124954 0 125010 800
rect 125506 0 125562 800
rect 126150 0 126206 800
rect 126702 0 126758 800
rect 127346 0 127402 800
rect 127990 0 128046 800
rect 128542 0 128598 800
rect 129186 0 129242 800
rect 129738 0 129794 800
rect 130382 0 130438 800
rect 131026 0 131082 800
rect 131578 0 131634 800
rect 132222 0 132278 800
rect 132866 0 132922 800
rect 133418 0 133474 800
rect 134062 0 134118 800
rect 134614 0 134670 800
rect 135258 0 135314 800
rect 135902 0 135958 800
rect 136454 0 136510 800
rect 137098 0 137154 800
rect 137650 0 137706 800
rect 138294 0 138350 800
rect 138938 0 138994 800
rect 139490 0 139546 800
rect 140134 0 140190 800
rect 140686 0 140742 800
rect 141330 0 141386 800
rect 141974 0 142030 800
rect 142526 0 142582 800
rect 143170 0 143226 800
rect 143814 0 143870 800
rect 144366 0 144422 800
rect 145010 0 145066 800
rect 145562 0 145618 800
rect 146206 0 146262 800
rect 146850 0 146906 800
rect 147402 0 147458 800
rect 148046 0 148102 800
rect 148598 0 148654 800
rect 149242 0 149298 800
rect 149886 0 149942 800
rect 150438 0 150494 800
rect 151082 0 151138 800
rect 151634 0 151690 800
rect 152278 0 152334 800
rect 152922 0 152978 800
rect 153474 0 153530 800
rect 154118 0 154174 800
rect 154670 0 154726 800
rect 155314 0 155370 800
rect 155958 0 156014 800
rect 156510 0 156566 800
rect 157154 0 157210 800
rect 157798 0 157854 800
rect 158350 0 158406 800
rect 158994 0 159050 800
rect 159546 0 159602 800
rect 160190 0 160246 800
rect 160834 0 160890 800
rect 161386 0 161442 800
rect 162030 0 162086 800
rect 162582 0 162638 800
rect 163226 0 163282 800
rect 163870 0 163926 800
rect 164422 0 164478 800
rect 165066 0 165122 800
rect 165618 0 165674 800
rect 166262 0 166318 800
rect 166906 0 166962 800
rect 167458 0 167514 800
rect 168102 0 168158 800
rect 168746 0 168802 800
rect 169298 0 169354 800
rect 169942 0 169998 800
rect 170494 0 170550 800
rect 171138 0 171194 800
rect 171782 0 171838 800
rect 172334 0 172390 800
rect 172978 0 173034 800
rect 173530 0 173586 800
rect 174174 0 174230 800
rect 174818 0 174874 800
rect 175370 0 175426 800
rect 176014 0 176070 800
rect 176566 0 176622 800
rect 177210 0 177266 800
rect 177854 0 177910 800
rect 178406 0 178462 800
rect 179050 0 179106 800
rect 179694 0 179750 800
rect 180246 0 180302 800
rect 180890 0 180946 800
rect 181442 0 181498 800
rect 182086 0 182142 800
rect 182730 0 182786 800
rect 183282 0 183338 800
rect 183926 0 183982 800
rect 184478 0 184534 800
rect 185122 0 185178 800
rect 185766 0 185822 800
rect 186318 0 186374 800
rect 186962 0 187018 800
rect 187514 0 187570 800
rect 188158 0 188214 800
rect 188802 0 188858 800
rect 189354 0 189410 800
rect 189998 0 190054 800
rect 190550 0 190606 800
rect 191194 0 191250 800
rect 191838 0 191894 800
rect 192390 0 192446 800
rect 193034 0 193090 800
rect 193678 0 193734 800
rect 194230 0 194286 800
rect 194874 0 194930 800
rect 195426 0 195482 800
rect 196070 0 196126 800
rect 196714 0 196770 800
rect 197266 0 197322 800
rect 197910 0 197966 800
rect 198462 0 198518 800
rect 199106 0 199162 800
rect 199750 0 199806 800
rect 200302 0 200358 800
rect 200946 0 201002 800
rect 201498 0 201554 800
rect 202142 0 202198 800
rect 202786 0 202842 800
rect 203338 0 203394 800
rect 203982 0 204038 800
rect 204626 0 204682 800
rect 205178 0 205234 800
rect 205822 0 205878 800
rect 206374 0 206430 800
rect 207018 0 207074 800
rect 207662 0 207718 800
rect 208214 0 208270 800
rect 208858 0 208914 800
rect 209410 0 209466 800
rect 210054 0 210110 800
rect 210698 0 210754 800
rect 211250 0 211306 800
rect 211894 0 211950 800
rect 212446 0 212502 800
rect 213090 0 213146 800
rect 213734 0 213790 800
rect 214286 0 214342 800
rect 214930 0 214986 800
rect 215574 0 215630 800
rect 216126 0 216182 800
rect 216770 0 216826 800
rect 217322 0 217378 800
rect 217966 0 218022 800
rect 218610 0 218666 800
rect 219162 0 219218 800
rect 219806 0 219862 800
rect 220358 0 220414 800
rect 221002 0 221058 800
rect 221646 0 221702 800
rect 222198 0 222254 800
rect 222842 0 222898 800
rect 223394 0 223450 800
rect 224038 0 224094 800
rect 224682 0 224738 800
rect 225234 0 225290 800
rect 225878 0 225934 800
rect 226430 0 226486 800
rect 227074 0 227130 800
rect 227718 0 227774 800
rect 228270 0 228326 800
rect 228914 0 228970 800
rect 229558 0 229614 800
rect 230110 0 230166 800
rect 230754 0 230810 800
rect 231306 0 231362 800
rect 231950 0 232006 800
rect 232594 0 232650 800
rect 233146 0 233202 800
rect 233790 0 233846 800
rect 234342 0 234398 800
rect 234986 0 235042 800
rect 235630 0 235686 800
rect 236182 0 236238 800
rect 236826 0 236882 800
rect 237378 0 237434 800
rect 238022 0 238078 800
rect 238666 0 238722 800
rect 239218 0 239274 800
rect 239862 0 239918 800
rect 240506 0 240562 800
rect 241058 0 241114 800
rect 241702 0 241758 800
rect 242254 0 242310 800
rect 242898 0 242954 800
rect 243542 0 243598 800
rect 244094 0 244150 800
rect 244738 0 244794 800
rect 245290 0 245346 800
rect 245934 0 245990 800
rect 246578 0 246634 800
rect 247130 0 247186 800
rect 247774 0 247830 800
rect 248326 0 248382 800
rect 248970 0 249026 800
rect 249614 0 249670 800
rect 250166 0 250222 800
rect 250810 0 250866 800
rect 251454 0 251510 800
rect 252006 0 252062 800
rect 252650 0 252706 800
rect 253202 0 253258 800
rect 253846 0 253902 800
rect 254490 0 254546 800
rect 255042 0 255098 800
rect 255686 0 255742 800
rect 256238 0 256294 800
rect 256882 0 256938 800
rect 257526 0 257582 800
rect 258078 0 258134 800
rect 258722 0 258778 800
rect 259274 0 259330 800
rect 259918 0 259974 800
rect 260562 0 260618 800
rect 261114 0 261170 800
rect 261758 0 261814 800
rect 262310 0 262366 800
rect 262954 0 263010 800
rect 263598 0 263654 800
rect 264150 0 264206 800
rect 264794 0 264850 800
rect 265438 0 265494 800
rect 265990 0 266046 800
rect 266634 0 266690 800
rect 267186 0 267242 800
rect 267830 0 267886 800
rect 268474 0 268530 800
rect 269026 0 269082 800
rect 269670 0 269726 800
rect 270222 0 270278 800
rect 270866 0 270922 800
rect 271510 0 271566 800
rect 272062 0 272118 800
rect 272706 0 272762 800
rect 273258 0 273314 800
rect 273902 0 273958 800
rect 274546 0 274602 800
rect 275098 0 275154 800
rect 275742 0 275798 800
rect 276386 0 276442 800
rect 276938 0 276994 800
rect 277582 0 277638 800
rect 278134 0 278190 800
rect 278778 0 278834 800
rect 279422 0 279478 800
rect 279974 0 280030 800
rect 280618 0 280674 800
rect 281170 0 281226 800
rect 281814 0 281870 800
rect 282458 0 282514 800
rect 283010 0 283066 800
rect 283654 0 283710 800
rect 284206 0 284262 800
rect 284850 0 284906 800
rect 285494 0 285550 800
rect 286046 0 286102 800
rect 286690 0 286746 800
rect 287334 0 287390 800
rect 287886 0 287942 800
rect 288530 0 288586 800
rect 289082 0 289138 800
rect 289726 0 289782 800
rect 290370 0 290426 800
rect 290922 0 290978 800
rect 291566 0 291622 800
rect 292118 0 292174 800
rect 292762 0 292818 800
rect 293406 0 293462 800
rect 293958 0 294014 800
rect 294602 0 294658 800
rect 295154 0 295210 800
rect 295798 0 295854 800
rect 296442 0 296498 800
rect 296994 0 297050 800
rect 297638 0 297694 800
<< obsm2 >>
rect 296 297144 1250 297200
rect 1418 297144 3826 297200
rect 3994 297144 6402 297200
rect 6570 297144 9070 297200
rect 9238 297144 11646 297200
rect 11814 297144 14314 297200
rect 14482 297144 16890 297200
rect 17058 297144 19466 297200
rect 19634 297144 22134 297200
rect 22302 297144 24710 297200
rect 24878 297144 27378 297200
rect 27546 297144 29954 297200
rect 30122 297144 32530 297200
rect 32698 297144 35198 297200
rect 35366 297144 37774 297200
rect 37942 297144 40442 297200
rect 40610 297144 43018 297200
rect 43186 297144 45686 297200
rect 45854 297144 48262 297200
rect 48430 297144 50838 297200
rect 51006 297144 53506 297200
rect 53674 297144 56082 297200
rect 56250 297144 58750 297200
rect 58918 297144 61326 297200
rect 61494 297144 63902 297200
rect 64070 297144 66570 297200
rect 66738 297144 69146 297200
rect 69314 297144 71814 297200
rect 71982 297144 74390 297200
rect 74558 297144 76966 297200
rect 77134 297144 79634 297200
rect 79802 297144 82210 297200
rect 82378 297144 84878 297200
rect 85046 297144 87454 297200
rect 87622 297144 90122 297200
rect 90290 297144 92698 297200
rect 92866 297144 95274 297200
rect 95442 297144 97942 297200
rect 98110 297144 100518 297200
rect 100686 297144 103186 297200
rect 103354 297144 105762 297200
rect 105930 297144 108338 297200
rect 108506 297144 111006 297200
rect 111174 297144 113582 297200
rect 113750 297144 116250 297200
rect 116418 297144 118826 297200
rect 118994 297144 121402 297200
rect 121570 297144 124070 297200
rect 124238 297144 126646 297200
rect 126814 297144 129314 297200
rect 129482 297144 131890 297200
rect 132058 297144 134558 297200
rect 134726 297144 137134 297200
rect 137302 297144 139710 297200
rect 139878 297144 142378 297200
rect 142546 297144 144954 297200
rect 145122 297144 147622 297200
rect 147790 297144 150198 297200
rect 150366 297144 152774 297200
rect 152942 297144 155442 297200
rect 155610 297144 158018 297200
rect 158186 297144 160686 297200
rect 160854 297144 163262 297200
rect 163430 297144 165838 297200
rect 166006 297144 168506 297200
rect 168674 297144 171082 297200
rect 171250 297144 173750 297200
rect 173918 297144 176326 297200
rect 176494 297144 178994 297200
rect 179162 297144 181570 297200
rect 181738 297144 184146 297200
rect 184314 297144 186814 297200
rect 186982 297144 189390 297200
rect 189558 297144 192058 297200
rect 192226 297144 194634 297200
rect 194802 297144 197210 297200
rect 197378 297144 199878 297200
rect 200046 297144 202454 297200
rect 202622 297144 205122 297200
rect 205290 297144 207698 297200
rect 207866 297144 210274 297200
rect 210442 297144 212942 297200
rect 213110 297144 215518 297200
rect 215686 297144 218186 297200
rect 218354 297144 220762 297200
rect 220930 297144 223430 297200
rect 223598 297144 226006 297200
rect 226174 297144 228582 297200
rect 228750 297144 231250 297200
rect 231418 297144 233826 297200
rect 233994 297144 236494 297200
rect 236662 297144 239070 297200
rect 239238 297144 241646 297200
rect 241814 297144 244314 297200
rect 244482 297144 246890 297200
rect 247058 297144 249558 297200
rect 249726 297144 252134 297200
rect 252302 297144 254710 297200
rect 254878 297144 257378 297200
rect 257546 297144 259954 297200
rect 260122 297144 262622 297200
rect 262790 297144 265198 297200
rect 265366 297144 267866 297200
rect 268034 297144 270442 297200
rect 270610 297144 273018 297200
rect 273186 297144 275686 297200
rect 275854 297144 278262 297200
rect 278430 297144 280930 297200
rect 281098 297144 283506 297200
rect 283674 297144 286082 297200
rect 286250 297144 288750 297200
rect 288918 297144 291326 297200
rect 291494 297144 293994 297200
rect 294162 297144 296570 297200
rect 296738 297144 297692 297200
rect 296 856 297692 297144
rect 406 800 790 856
rect 958 800 1434 856
rect 1602 800 1986 856
rect 2154 800 2630 856
rect 2798 800 3274 856
rect 3442 800 3826 856
rect 3994 800 4470 856
rect 4638 800 5022 856
rect 5190 800 5666 856
rect 5834 800 6310 856
rect 6478 800 6862 856
rect 7030 800 7506 856
rect 7674 800 8058 856
rect 8226 800 8702 856
rect 8870 800 9346 856
rect 9514 800 9898 856
rect 10066 800 10542 856
rect 10710 800 11094 856
rect 11262 800 11738 856
rect 11906 800 12382 856
rect 12550 800 12934 856
rect 13102 800 13578 856
rect 13746 800 14222 856
rect 14390 800 14774 856
rect 14942 800 15418 856
rect 15586 800 15970 856
rect 16138 800 16614 856
rect 16782 800 17258 856
rect 17426 800 17810 856
rect 17978 800 18454 856
rect 18622 800 19006 856
rect 19174 800 19650 856
rect 19818 800 20294 856
rect 20462 800 20846 856
rect 21014 800 21490 856
rect 21658 800 22042 856
rect 22210 800 22686 856
rect 22854 800 23330 856
rect 23498 800 23882 856
rect 24050 800 24526 856
rect 24694 800 25170 856
rect 25338 800 25722 856
rect 25890 800 26366 856
rect 26534 800 26918 856
rect 27086 800 27562 856
rect 27730 800 28206 856
rect 28374 800 28758 856
rect 28926 800 29402 856
rect 29570 800 29954 856
rect 30122 800 30598 856
rect 30766 800 31242 856
rect 31410 800 31794 856
rect 31962 800 32438 856
rect 32606 800 32990 856
rect 33158 800 33634 856
rect 33802 800 34278 856
rect 34446 800 34830 856
rect 34998 800 35474 856
rect 35642 800 36118 856
rect 36286 800 36670 856
rect 36838 800 37314 856
rect 37482 800 37866 856
rect 38034 800 38510 856
rect 38678 800 39154 856
rect 39322 800 39706 856
rect 39874 800 40350 856
rect 40518 800 40902 856
rect 41070 800 41546 856
rect 41714 800 42190 856
rect 42358 800 42742 856
rect 42910 800 43386 856
rect 43554 800 43938 856
rect 44106 800 44582 856
rect 44750 800 45226 856
rect 45394 800 45778 856
rect 45946 800 46422 856
rect 46590 800 46974 856
rect 47142 800 47618 856
rect 47786 800 48262 856
rect 48430 800 48814 856
rect 48982 800 49458 856
rect 49626 800 50102 856
rect 50270 800 50654 856
rect 50822 800 51298 856
rect 51466 800 51850 856
rect 52018 800 52494 856
rect 52662 800 53138 856
rect 53306 800 53690 856
rect 53858 800 54334 856
rect 54502 800 54886 856
rect 55054 800 55530 856
rect 55698 800 56174 856
rect 56342 800 56726 856
rect 56894 800 57370 856
rect 57538 800 57922 856
rect 58090 800 58566 856
rect 58734 800 59210 856
rect 59378 800 59762 856
rect 59930 800 60406 856
rect 60574 800 61050 856
rect 61218 800 61602 856
rect 61770 800 62246 856
rect 62414 800 62798 856
rect 62966 800 63442 856
rect 63610 800 64086 856
rect 64254 800 64638 856
rect 64806 800 65282 856
rect 65450 800 65834 856
rect 66002 800 66478 856
rect 66646 800 67122 856
rect 67290 800 67674 856
rect 67842 800 68318 856
rect 68486 800 68870 856
rect 69038 800 69514 856
rect 69682 800 70158 856
rect 70326 800 70710 856
rect 70878 800 71354 856
rect 71522 800 71998 856
rect 72166 800 72550 856
rect 72718 800 73194 856
rect 73362 800 73746 856
rect 73914 800 74390 856
rect 74558 800 75034 856
rect 75202 800 75586 856
rect 75754 800 76230 856
rect 76398 800 76782 856
rect 76950 800 77426 856
rect 77594 800 78070 856
rect 78238 800 78622 856
rect 78790 800 79266 856
rect 79434 800 79818 856
rect 79986 800 80462 856
rect 80630 800 81106 856
rect 81274 800 81658 856
rect 81826 800 82302 856
rect 82470 800 82854 856
rect 83022 800 83498 856
rect 83666 800 84142 856
rect 84310 800 84694 856
rect 84862 800 85338 856
rect 85506 800 85982 856
rect 86150 800 86534 856
rect 86702 800 87178 856
rect 87346 800 87730 856
rect 87898 800 88374 856
rect 88542 800 89018 856
rect 89186 800 89570 856
rect 89738 800 90214 856
rect 90382 800 90766 856
rect 90934 800 91410 856
rect 91578 800 92054 856
rect 92222 800 92606 856
rect 92774 800 93250 856
rect 93418 800 93802 856
rect 93970 800 94446 856
rect 94614 800 95090 856
rect 95258 800 95642 856
rect 95810 800 96286 856
rect 96454 800 96930 856
rect 97098 800 97482 856
rect 97650 800 98126 856
rect 98294 800 98678 856
rect 98846 800 99322 856
rect 99490 800 99966 856
rect 100134 800 100518 856
rect 100686 800 101162 856
rect 101330 800 101714 856
rect 101882 800 102358 856
rect 102526 800 103002 856
rect 103170 800 103554 856
rect 103722 800 104198 856
rect 104366 800 104750 856
rect 104918 800 105394 856
rect 105562 800 106038 856
rect 106206 800 106590 856
rect 106758 800 107234 856
rect 107402 800 107878 856
rect 108046 800 108430 856
rect 108598 800 109074 856
rect 109242 800 109626 856
rect 109794 800 110270 856
rect 110438 800 110914 856
rect 111082 800 111466 856
rect 111634 800 112110 856
rect 112278 800 112662 856
rect 112830 800 113306 856
rect 113474 800 113950 856
rect 114118 800 114502 856
rect 114670 800 115146 856
rect 115314 800 115698 856
rect 115866 800 116342 856
rect 116510 800 116986 856
rect 117154 800 117538 856
rect 117706 800 118182 856
rect 118350 800 118734 856
rect 118902 800 119378 856
rect 119546 800 120022 856
rect 120190 800 120574 856
rect 120742 800 121218 856
rect 121386 800 121862 856
rect 122030 800 122414 856
rect 122582 800 123058 856
rect 123226 800 123610 856
rect 123778 800 124254 856
rect 124422 800 124898 856
rect 125066 800 125450 856
rect 125618 800 126094 856
rect 126262 800 126646 856
rect 126814 800 127290 856
rect 127458 800 127934 856
rect 128102 800 128486 856
rect 128654 800 129130 856
rect 129298 800 129682 856
rect 129850 800 130326 856
rect 130494 800 130970 856
rect 131138 800 131522 856
rect 131690 800 132166 856
rect 132334 800 132810 856
rect 132978 800 133362 856
rect 133530 800 134006 856
rect 134174 800 134558 856
rect 134726 800 135202 856
rect 135370 800 135846 856
rect 136014 800 136398 856
rect 136566 800 137042 856
rect 137210 800 137594 856
rect 137762 800 138238 856
rect 138406 800 138882 856
rect 139050 800 139434 856
rect 139602 800 140078 856
rect 140246 800 140630 856
rect 140798 800 141274 856
rect 141442 800 141918 856
rect 142086 800 142470 856
rect 142638 800 143114 856
rect 143282 800 143758 856
rect 143926 800 144310 856
rect 144478 800 144954 856
rect 145122 800 145506 856
rect 145674 800 146150 856
rect 146318 800 146794 856
rect 146962 800 147346 856
rect 147514 800 147990 856
rect 148158 800 148542 856
rect 148710 800 149186 856
rect 149354 800 149830 856
rect 149998 800 150382 856
rect 150550 800 151026 856
rect 151194 800 151578 856
rect 151746 800 152222 856
rect 152390 800 152866 856
rect 153034 800 153418 856
rect 153586 800 154062 856
rect 154230 800 154614 856
rect 154782 800 155258 856
rect 155426 800 155902 856
rect 156070 800 156454 856
rect 156622 800 157098 856
rect 157266 800 157742 856
rect 157910 800 158294 856
rect 158462 800 158938 856
rect 159106 800 159490 856
rect 159658 800 160134 856
rect 160302 800 160778 856
rect 160946 800 161330 856
rect 161498 800 161974 856
rect 162142 800 162526 856
rect 162694 800 163170 856
rect 163338 800 163814 856
rect 163982 800 164366 856
rect 164534 800 165010 856
rect 165178 800 165562 856
rect 165730 800 166206 856
rect 166374 800 166850 856
rect 167018 800 167402 856
rect 167570 800 168046 856
rect 168214 800 168690 856
rect 168858 800 169242 856
rect 169410 800 169886 856
rect 170054 800 170438 856
rect 170606 800 171082 856
rect 171250 800 171726 856
rect 171894 800 172278 856
rect 172446 800 172922 856
rect 173090 800 173474 856
rect 173642 800 174118 856
rect 174286 800 174762 856
rect 174930 800 175314 856
rect 175482 800 175958 856
rect 176126 800 176510 856
rect 176678 800 177154 856
rect 177322 800 177798 856
rect 177966 800 178350 856
rect 178518 800 178994 856
rect 179162 800 179638 856
rect 179806 800 180190 856
rect 180358 800 180834 856
rect 181002 800 181386 856
rect 181554 800 182030 856
rect 182198 800 182674 856
rect 182842 800 183226 856
rect 183394 800 183870 856
rect 184038 800 184422 856
rect 184590 800 185066 856
rect 185234 800 185710 856
rect 185878 800 186262 856
rect 186430 800 186906 856
rect 187074 800 187458 856
rect 187626 800 188102 856
rect 188270 800 188746 856
rect 188914 800 189298 856
rect 189466 800 189942 856
rect 190110 800 190494 856
rect 190662 800 191138 856
rect 191306 800 191782 856
rect 191950 800 192334 856
rect 192502 800 192978 856
rect 193146 800 193622 856
rect 193790 800 194174 856
rect 194342 800 194818 856
rect 194986 800 195370 856
rect 195538 800 196014 856
rect 196182 800 196658 856
rect 196826 800 197210 856
rect 197378 800 197854 856
rect 198022 800 198406 856
rect 198574 800 199050 856
rect 199218 800 199694 856
rect 199862 800 200246 856
rect 200414 800 200890 856
rect 201058 800 201442 856
rect 201610 800 202086 856
rect 202254 800 202730 856
rect 202898 800 203282 856
rect 203450 800 203926 856
rect 204094 800 204570 856
rect 204738 800 205122 856
rect 205290 800 205766 856
rect 205934 800 206318 856
rect 206486 800 206962 856
rect 207130 800 207606 856
rect 207774 800 208158 856
rect 208326 800 208802 856
rect 208970 800 209354 856
rect 209522 800 209998 856
rect 210166 800 210642 856
rect 210810 800 211194 856
rect 211362 800 211838 856
rect 212006 800 212390 856
rect 212558 800 213034 856
rect 213202 800 213678 856
rect 213846 800 214230 856
rect 214398 800 214874 856
rect 215042 800 215518 856
rect 215686 800 216070 856
rect 216238 800 216714 856
rect 216882 800 217266 856
rect 217434 800 217910 856
rect 218078 800 218554 856
rect 218722 800 219106 856
rect 219274 800 219750 856
rect 219918 800 220302 856
rect 220470 800 220946 856
rect 221114 800 221590 856
rect 221758 800 222142 856
rect 222310 800 222786 856
rect 222954 800 223338 856
rect 223506 800 223982 856
rect 224150 800 224626 856
rect 224794 800 225178 856
rect 225346 800 225822 856
rect 225990 800 226374 856
rect 226542 800 227018 856
rect 227186 800 227662 856
rect 227830 800 228214 856
rect 228382 800 228858 856
rect 229026 800 229502 856
rect 229670 800 230054 856
rect 230222 800 230698 856
rect 230866 800 231250 856
rect 231418 800 231894 856
rect 232062 800 232538 856
rect 232706 800 233090 856
rect 233258 800 233734 856
rect 233902 800 234286 856
rect 234454 800 234930 856
rect 235098 800 235574 856
rect 235742 800 236126 856
rect 236294 800 236770 856
rect 236938 800 237322 856
rect 237490 800 237966 856
rect 238134 800 238610 856
rect 238778 800 239162 856
rect 239330 800 239806 856
rect 239974 800 240450 856
rect 240618 800 241002 856
rect 241170 800 241646 856
rect 241814 800 242198 856
rect 242366 800 242842 856
rect 243010 800 243486 856
rect 243654 800 244038 856
rect 244206 800 244682 856
rect 244850 800 245234 856
rect 245402 800 245878 856
rect 246046 800 246522 856
rect 246690 800 247074 856
rect 247242 800 247718 856
rect 247886 800 248270 856
rect 248438 800 248914 856
rect 249082 800 249558 856
rect 249726 800 250110 856
rect 250278 800 250754 856
rect 250922 800 251398 856
rect 251566 800 251950 856
rect 252118 800 252594 856
rect 252762 800 253146 856
rect 253314 800 253790 856
rect 253958 800 254434 856
rect 254602 800 254986 856
rect 255154 800 255630 856
rect 255798 800 256182 856
rect 256350 800 256826 856
rect 256994 800 257470 856
rect 257638 800 258022 856
rect 258190 800 258666 856
rect 258834 800 259218 856
rect 259386 800 259862 856
rect 260030 800 260506 856
rect 260674 800 261058 856
rect 261226 800 261702 856
rect 261870 800 262254 856
rect 262422 800 262898 856
rect 263066 800 263542 856
rect 263710 800 264094 856
rect 264262 800 264738 856
rect 264906 800 265382 856
rect 265550 800 265934 856
rect 266102 800 266578 856
rect 266746 800 267130 856
rect 267298 800 267774 856
rect 267942 800 268418 856
rect 268586 800 268970 856
rect 269138 800 269614 856
rect 269782 800 270166 856
rect 270334 800 270810 856
rect 270978 800 271454 856
rect 271622 800 272006 856
rect 272174 800 272650 856
rect 272818 800 273202 856
rect 273370 800 273846 856
rect 274014 800 274490 856
rect 274658 800 275042 856
rect 275210 800 275686 856
rect 275854 800 276330 856
rect 276498 800 276882 856
rect 277050 800 277526 856
rect 277694 800 278078 856
rect 278246 800 278722 856
rect 278890 800 279366 856
rect 279534 800 279918 856
rect 280086 800 280562 856
rect 280730 800 281114 856
rect 281282 800 281758 856
rect 281926 800 282402 856
rect 282570 800 282954 856
rect 283122 800 283598 856
rect 283766 800 284150 856
rect 284318 800 284794 856
rect 284962 800 285438 856
rect 285606 800 285990 856
rect 286158 800 286634 856
rect 286802 800 287278 856
rect 287446 800 287830 856
rect 287998 800 288474 856
rect 288642 800 289026 856
rect 289194 800 289670 856
rect 289838 800 290314 856
rect 290482 800 290866 856
rect 291034 800 291510 856
rect 291678 800 292062 856
rect 292230 800 292706 856
rect 292874 800 293350 856
rect 293518 800 293902 856
rect 294070 800 294546 856
rect 294714 800 295098 856
rect 295266 800 295742 856
rect 295910 800 296386 856
rect 296554 800 296938 856
rect 297106 800 297582 856
<< metal3 >>
rect 297200 248208 298000 248328
rect 0 148928 800 149048
rect 297200 148928 298000 149048
rect 297200 49648 298000 49768
<< obsm3 >>
rect 800 248408 297200 295425
rect 800 248128 297120 248408
rect 800 149128 297200 248128
rect 880 148848 297120 149128
rect 800 49848 297200 148848
rect 800 49568 297120 49848
rect 800 2143 297200 49568
<< metal4 >>
rect 4208 2128 4528 295440
rect 4868 2176 5188 295392
rect 5528 2176 5848 295392
rect 6188 2176 6508 295392
rect 19568 2128 19888 295440
rect 20228 2176 20548 295392
rect 20888 2176 21208 295392
rect 21548 2176 21868 295392
rect 34928 2128 35248 295440
rect 35588 2176 35908 295392
rect 36248 2176 36568 295392
rect 36908 2176 37228 295392
rect 50288 2128 50608 295440
rect 50948 2176 51268 295392
rect 51608 2176 51928 295392
rect 52268 2176 52588 295392
rect 65648 2128 65968 295440
rect 66308 2176 66628 295392
rect 66968 2176 67288 295392
rect 67628 2176 67948 295392
rect 81008 2128 81328 295440
rect 81668 2176 81988 295392
rect 82328 2176 82648 295392
rect 82988 2176 83308 295392
rect 96368 2128 96688 295440
rect 97028 2176 97348 295392
rect 97688 2176 98008 295392
rect 98348 2176 98668 295392
rect 111728 2128 112048 295440
rect 112388 2176 112708 295392
rect 113048 2176 113368 295392
rect 113708 2176 114028 295392
rect 127088 2128 127408 295440
rect 127748 2176 128068 295392
rect 128408 2176 128728 295392
rect 129068 2176 129388 295392
rect 142448 2128 142768 295440
rect 143108 2176 143428 295392
rect 143768 2176 144088 295392
rect 144428 2176 144748 295392
rect 157808 2128 158128 295440
rect 158468 2176 158788 295392
rect 159128 2176 159448 295392
rect 159788 2176 160108 295392
rect 173168 2128 173488 295440
rect 173828 2176 174148 295392
rect 174488 2176 174808 295392
rect 175148 2176 175468 295392
rect 188528 2128 188848 295440
rect 189188 2176 189508 295392
rect 189848 2176 190168 295392
rect 190508 2176 190828 295392
rect 203888 2128 204208 295440
rect 204548 2176 204868 295392
rect 205208 2176 205528 295392
rect 205868 2176 206188 295392
rect 219248 2128 219568 295440
rect 219908 2176 220228 295392
rect 220568 2176 220888 295392
rect 221228 2176 221548 295392
rect 234608 2128 234928 295440
rect 235268 2176 235588 295392
rect 235928 2176 236248 295392
rect 236588 2176 236908 295392
rect 249968 2128 250288 295440
rect 250628 2176 250948 295392
rect 251288 2176 251608 295392
rect 251948 2176 252268 295392
rect 265328 2128 265648 295440
rect 265988 2176 266308 295392
rect 266648 2176 266968 295392
rect 267308 2176 267628 295392
rect 280688 2128 281008 295440
rect 281348 2176 281668 295392
rect 282008 2176 282328 295392
rect 282668 2176 282988 295392
rect 296048 2128 296368 295440
<< obsm4 >>
rect 2451 2619 4128 292773
rect 4608 2619 4788 292773
rect 5268 2619 5448 292773
rect 5928 2619 6108 292773
rect 6588 2619 19488 292773
rect 19968 2619 20148 292773
rect 20628 2619 20808 292773
rect 21288 2619 21468 292773
rect 21948 2619 34848 292773
rect 35328 2619 35508 292773
rect 35988 2619 36168 292773
rect 36648 2619 36828 292773
rect 37308 2619 50208 292773
rect 50688 2619 50868 292773
rect 51348 2619 51528 292773
rect 52008 2619 52188 292773
rect 52668 2619 65568 292773
rect 66048 2619 66228 292773
rect 66708 2619 66888 292773
rect 67368 2619 67548 292773
rect 68028 2619 80928 292773
rect 81408 2619 81588 292773
rect 82068 2619 82248 292773
rect 82728 2619 82908 292773
rect 83388 2619 96288 292773
rect 96768 2619 96948 292773
rect 97428 2619 97608 292773
rect 98088 2619 98268 292773
rect 98748 2619 111648 292773
rect 112128 2619 112308 292773
rect 112788 2619 112968 292773
rect 113448 2619 113628 292773
rect 114108 2619 127008 292773
rect 127488 2619 127668 292773
rect 128148 2619 128328 292773
rect 128808 2619 128988 292773
rect 129468 2619 142368 292773
rect 142848 2619 143028 292773
rect 143508 2619 143688 292773
rect 144168 2619 144348 292773
rect 144828 2619 157728 292773
rect 158208 2619 158388 292773
rect 158868 2619 159048 292773
rect 159528 2619 159708 292773
rect 160188 2619 173088 292773
rect 173568 2619 173748 292773
rect 174228 2619 174408 292773
rect 174888 2619 175068 292773
rect 175548 2619 188448 292773
rect 188928 2619 189108 292773
rect 189588 2619 189768 292773
rect 190248 2619 190428 292773
rect 190908 2619 203808 292773
rect 204288 2619 204468 292773
rect 204948 2619 205128 292773
rect 205608 2619 205788 292773
rect 206268 2619 219168 292773
rect 219648 2619 219828 292773
rect 220308 2619 220488 292773
rect 220968 2619 221148 292773
rect 221628 2619 234528 292773
rect 235008 2619 235188 292773
rect 235668 2619 235848 292773
rect 236328 2619 236508 292773
rect 236988 2619 249888 292773
rect 250368 2619 250548 292773
rect 251028 2619 251208 292773
rect 251688 2619 251868 292773
rect 252348 2619 265248 292773
rect 265728 2619 265908 292773
rect 266388 2619 266568 292773
rect 267048 2619 267228 292773
rect 267708 2619 280608 292773
rect 281088 2619 281268 292773
rect 281748 2619 281928 292773
rect 282408 2619 282588 292773
rect 283068 2619 290661 292773
<< labels >>
rlabel metal2 s 1306 297200 1362 298000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 79690 297200 79746 298000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 87510 297200 87566 298000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 95330 297200 95386 298000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 103242 297200 103298 298000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 111062 297200 111118 298000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 118882 297200 118938 298000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 126702 297200 126758 298000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 134614 297200 134670 298000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 142434 297200 142490 298000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 150254 297200 150310 298000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 9126 297200 9182 298000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 158074 297200 158130 298000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 165894 297200 165950 298000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 173806 297200 173862 298000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 181626 297200 181682 298000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 189446 297200 189502 298000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 197266 297200 197322 298000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 205178 297200 205234 298000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 212998 297200 213054 298000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 220818 297200 220874 298000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 228638 297200 228694 298000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 16946 297200 17002 298000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 236550 297200 236606 298000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 244370 297200 244426 298000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 252190 297200 252246 298000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 260010 297200 260066 298000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 267922 297200 267978 298000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 275742 297200 275798 298000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 283562 297200 283618 298000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 291382 297200 291438 298000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 24766 297200 24822 298000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 32586 297200 32642 298000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 40498 297200 40554 298000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 48318 297200 48374 298000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 56138 297200 56194 298000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 63958 297200 64014 298000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 71870 297200 71926 298000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3882 297200 3938 298000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 82266 297200 82322 298000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 90178 297200 90234 298000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 97998 297200 98054 298000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 105818 297200 105874 298000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 113638 297200 113694 298000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 121458 297200 121514 298000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 129370 297200 129426 298000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 137190 297200 137246 298000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 145010 297200 145066 298000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 152830 297200 152886 298000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 11702 297200 11758 298000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 160742 297200 160798 298000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 168562 297200 168618 298000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 176382 297200 176438 298000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 184202 297200 184258 298000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 192114 297200 192170 298000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 199934 297200 199990 298000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 207754 297200 207810 298000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 215574 297200 215630 298000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 223486 297200 223542 298000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 231306 297200 231362 298000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 19522 297200 19578 298000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 239126 297200 239182 298000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 246946 297200 247002 298000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 254766 297200 254822 298000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 262678 297200 262734 298000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 270498 297200 270554 298000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 278318 297200 278374 298000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 286138 297200 286194 298000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 294050 297200 294106 298000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 27434 297200 27490 298000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 35254 297200 35310 298000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 43074 297200 43130 298000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 50894 297200 50950 298000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 58806 297200 58862 298000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 66626 297200 66682 298000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 74446 297200 74502 298000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 6458 297200 6514 298000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 84934 297200 84990 298000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 92754 297200 92810 298000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 100574 297200 100630 298000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 108394 297200 108450 298000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 116306 297200 116362 298000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 124126 297200 124182 298000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 131946 297200 132002 298000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 139766 297200 139822 298000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 147678 297200 147734 298000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 155498 297200 155554 298000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 14370 297200 14426 298000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 163318 297200 163374 298000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 171138 297200 171194 298000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 179050 297200 179106 298000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 186870 297200 186926 298000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 194690 297200 194746 298000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 202510 297200 202566 298000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 210330 297200 210386 298000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 218242 297200 218298 298000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 226062 297200 226118 298000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 233882 297200 233938 298000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 22190 297200 22246 298000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 241702 297200 241758 298000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 249614 297200 249670 298000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 257434 297200 257490 298000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 265254 297200 265310 298000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 273074 297200 273130 298000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 280986 297200 281042 298000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 288806 297200 288862 298000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 296626 297200 296682 298000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 30010 297200 30066 298000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 37830 297200 37886 298000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 45742 297200 45798 298000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 53562 297200 53618 298000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 61382 297200 61438 298000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 69202 297200 69258 298000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 77022 297200 77078 298000 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 297200 148928 298000 149048 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 0 148928 800 149048 6 irq[1]
port 116 nsew signal output
rlabel metal3 s 297200 248208 298000 248328 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 247130 0 247186 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 248970 0 249026 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 250810 0 250866 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 252650 0 252706 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 254490 0 254546 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 256238 0 256294 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 258078 0 258134 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 259918 0 259974 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 261758 0 261814 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 263598 0 263654 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 265438 0 265494 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 267186 0 267242 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 269026 0 269082 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 270866 0 270922 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 272706 0 272762 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 274546 0 274602 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 276386 0 276442 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 278134 0 278190 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 279974 0 280030 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 281814 0 281870 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 283654 0 283710 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 285494 0 285550 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 287334 0 287390 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 289082 0 289138 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 290922 0 290978 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 292762 0 292818 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 294602 0 294658 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 296442 0 296498 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 106646 0 106702 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 119434 0 119490 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 126702 0 126758 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 148598 0 148654 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 150438 0 150494 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 152278 0 152334 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 154118 0 154174 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 155958 0 156014 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 159546 0 159602 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 161386 0 161442 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 163226 0 163282 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 166906 0 166962 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 170494 0 170550 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 172334 0 172390 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 174174 0 174230 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 176014 0 176070 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 177854 0 177910 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 179694 0 179750 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 181442 0 181498 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 183282 0 183338 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 185122 0 185178 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 186962 0 187018 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 188802 0 188858 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 190550 0 190606 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 192390 0 192446 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 194230 0 194286 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 196070 0 196126 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 197910 0 197966 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 199750 0 199806 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 201498 0 201554 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 203338 0 203394 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 205178 0 205234 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 207018 0 207074 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 208858 0 208914 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 210698 0 210754 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 212446 0 212502 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 214286 0 214342 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 216126 0 216182 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 217966 0 218022 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 219806 0 219862 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 221646 0 221702 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 223394 0 223450 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 225234 0 225290 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 227074 0 227130 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 228914 0 228970 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 230754 0 230810 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 232594 0 232650 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 234342 0 234398 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 236182 0 236238 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 238022 0 238078 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 239862 0 239918 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 241702 0 241758 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 243542 0 243598 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 245290 0 245346 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 247774 0 247830 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 249614 0 249670 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 251454 0 251510 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 253202 0 253258 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 255042 0 255098 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 256882 0 256938 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 258722 0 258778 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 260562 0 260618 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 262310 0 262366 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 264150 0 264206 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 83554 0 83610 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 265990 0 266046 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 267830 0 267886 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 269670 0 269726 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 271510 0 271566 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 273258 0 273314 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 275098 0 275154 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 276938 0 276994 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 278778 0 278834 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 280618 0 280674 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 282458 0 282514 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 85394 0 85450 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 284206 0 284262 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 286046 0 286102 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 287886 0 287942 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 289726 0 289782 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 291566 0 291622 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 293406 0 293462 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 295154 0 295210 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 296994 0 297050 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 89074 0 89130 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 92662 0 92718 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 94502 0 94558 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 96342 0 96398 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 98182 0 98238 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 100022 0 100078 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 103610 0 103666 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 105450 0 105506 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 107290 0 107346 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 109130 0 109186 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 110970 0 111026 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 114558 0 114614 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 116398 0 116454 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 118238 0 118294 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 120078 0 120134 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 125506 0 125562 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 127346 0 127402 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 129186 0 129242 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 131026 0 131082 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 132866 0 132922 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 136454 0 136510 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 138294 0 138350 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 140134 0 140190 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 141974 0 142030 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 143814 0 143870 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 145562 0 145618 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 147402 0 147458 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 149242 0 149298 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 151082 0 151138 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 152922 0 152978 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 154670 0 154726 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 72606 0 72662 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 156510 0 156566 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 158350 0 158406 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 160190 0 160246 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 162030 0 162086 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 165618 0 165674 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 167458 0 167514 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 169298 0 169354 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 171138 0 171194 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 172978 0 173034 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 174818 0 174874 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 176566 0 176622 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 178406 0 178462 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 180246 0 180302 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 182086 0 182142 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 183926 0 183982 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 185766 0 185822 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 187514 0 187570 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 189354 0 189410 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 191194 0 191250 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 76286 0 76342 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 193034 0 193090 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 194874 0 194930 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 196714 0 196770 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 198462 0 198518 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 200302 0 200358 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 202142 0 202198 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 203982 0 204038 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 205822 0 205878 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 207662 0 207718 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 209410 0 209466 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 211250 0 211306 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 213090 0 213146 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 214930 0 214986 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 216770 0 216826 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 218610 0 218666 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 220358 0 220414 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 222198 0 222254 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 224038 0 224094 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 225878 0 225934 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 227718 0 227774 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 229558 0 229614 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 231306 0 231362 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 233146 0 233202 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 234986 0 235042 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 236826 0 236882 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 238666 0 238722 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 240506 0 240562 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 242254 0 242310 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 244094 0 244150 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 245934 0 245990 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 81714 0 81770 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 248326 0 248382 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 250166 0 250222 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 252006 0 252062 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 253846 0 253902 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 255686 0 255742 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 257526 0 257582 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 259274 0 259330 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 261114 0 261170 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 262954 0 263010 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 264794 0 264850 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 266634 0 266690 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 268474 0 268530 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 270222 0 270278 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 272062 0 272118 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 273902 0 273958 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 275742 0 275798 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 277582 0 277638 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 279422 0 279478 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 281170 0 281226 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 283010 0 283066 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 284850 0 284906 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 286690 0 286746 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 288530 0 288586 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 290370 0 290426 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 292118 0 292174 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 293958 0 294014 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 295798 0 295854 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 297638 0 297694 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 109682 0 109738 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 122470 0 122526 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 126150 0 126206 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 140686 0 140742 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 144366 0 144422 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 148046 0 148102 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 149886 0 149942 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 151634 0 151690 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 153474 0 153530 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 155314 0 155370 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 158994 0 159050 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 160834 0 160890 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 162582 0 162638 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 164422 0 164478 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 166262 0 166318 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 168102 0 168158 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 169942 0 169998 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 175370 0 175426 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 177210 0 177266 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 180890 0 180946 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 182730 0 182786 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 184478 0 184534 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 186318 0 186374 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 188158 0 188214 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 191838 0 191894 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 193678 0 193734 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 195426 0 195482 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 197266 0 197322 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 199106 0 199162 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 200946 0 201002 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 202786 0 202842 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 204626 0 204682 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 206374 0 206430 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 208214 0 208270 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 210054 0 210110 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 211894 0 211950 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 213734 0 213790 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 215574 0 215630 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 217322 0 217378 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 219162 0 219218 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 221002 0 221058 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 222842 0 222898 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 224682 0 224738 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 226430 0 226486 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 228270 0 228326 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 230110 0 230166 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 231950 0 232006 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 233790 0 233846 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 235630 0 235686 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 237378 0 237434 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 239218 0 239274 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 241058 0 241114 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 242898 0 242954 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 244738 0 244794 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 246578 0 246634 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal3 s 297200 49648 298000 49768 6 user_clk
port 502 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 503 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 504 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_ack_o
port 505 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 wbs_adr_i[0]
port 506 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[10]
port 507 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_adr_i[11]
port 508 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wbs_adr_i[12]
port 509 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_adr_i[13]
port 510 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_adr_i[14]
port 511 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_adr_i[15]
port 512 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wbs_adr_i[16]
port 513 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 wbs_adr_i[17]
port 514 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 wbs_adr_i[18]
port 515 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 wbs_adr_i[19]
port 516 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_adr_i[1]
port 517 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 wbs_adr_i[20]
port 518 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 wbs_adr_i[21]
port 519 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wbs_adr_i[22]
port 520 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_adr_i[23]
port 521 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 wbs_adr_i[24]
port 522 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 wbs_adr_i[25]
port 523 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 wbs_adr_i[26]
port 524 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 wbs_adr_i[27]
port 525 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 wbs_adr_i[28]
port 526 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 wbs_adr_i[29]
port 527 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[2]
port 528 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 wbs_adr_i[30]
port 529 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 wbs_adr_i[31]
port 530 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_adr_i[3]
port 531 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_adr_i[4]
port 532 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_adr_i[5]
port 533 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_adr_i[6]
port 534 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_adr_i[7]
port 535 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[8]
port 536 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_adr_i[9]
port 537 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_cyc_i
port 538 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_dat_i[0]
port 539 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_i[10]
port 540 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_i[11]
port 541 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_i[12]
port 542 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 wbs_dat_i[13]
port 543 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_dat_i[14]
port 544 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_i[15]
port 545 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 wbs_dat_i[16]
port 546 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 wbs_dat_i[17]
port 547 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 wbs_dat_i[18]
port 548 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_i[19]
port 549 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_i[1]
port 550 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 wbs_dat_i[20]
port 551 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 wbs_dat_i[21]
port 552 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 wbs_dat_i[22]
port 553 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 wbs_dat_i[23]
port 554 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 wbs_dat_i[24]
port 555 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 wbs_dat_i[25]
port 556 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wbs_dat_i[26]
port 557 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 wbs_dat_i[27]
port 558 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 wbs_dat_i[28]
port 559 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 wbs_dat_i[29]
port 560 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_i[2]
port 561 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 wbs_dat_i[30]
port 562 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 wbs_dat_i[31]
port 563 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_i[3]
port 564 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_i[4]
port 565 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_dat_i[5]
port 566 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_dat_i[6]
port 567 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_i[7]
port 568 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_i[8]
port 569 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_i[9]
port 570 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_o[0]
port 571 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_o[10]
port 572 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_o[11]
port 573 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_o[12]
port 574 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 wbs_dat_o[13]
port 575 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 wbs_dat_o[14]
port 576 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_o[15]
port 577 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 wbs_dat_o[16]
port 578 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 wbs_dat_o[17]
port 579 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 wbs_dat_o[18]
port 580 nsew signal output
rlabel metal2 s 42246 0 42302 800 6 wbs_dat_o[19]
port 581 nsew signal output
rlabel metal2 s 7562 0 7618 800 6 wbs_dat_o[1]
port 582 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 wbs_dat_o[20]
port 583 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 wbs_dat_o[21]
port 584 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 wbs_dat_o[22]
port 585 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 wbs_dat_o[23]
port 586 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 wbs_dat_o[24]
port 587 nsew signal output
rlabel metal2 s 53194 0 53250 800 6 wbs_dat_o[25]
port 588 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 wbs_dat_o[26]
port 589 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 wbs_dat_o[27]
port 590 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 wbs_dat_o[28]
port 591 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 wbs_dat_o[29]
port 592 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[2]
port 593 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 wbs_dat_o[30]
port 594 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 wbs_dat_o[31]
port 595 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_o[3]
port 596 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[4]
port 597 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_o[5]
port 598 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_o[6]
port 599 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_o[7]
port 600 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_o[8]
port 601 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_o[9]
port 602 nsew signal output
rlabel metal2 s 5722 0 5778 800 6 wbs_sel_i[0]
port 603 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_sel_i[1]
port 604 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_sel_i[2]
port 605 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_sel_i[3]
port 606 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_stb_i
port 607 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_we_i
port 608 nsew signal input
rlabel metal4 s 280688 2128 281008 295440 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 295440 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 295440 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 295440 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 295440 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 295440 6 vccd1
port 614 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 295440 6 vccd1
port 615 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 295440 6 vccd1
port 616 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 295440 6 vccd1
port 617 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 295440 6 vccd1
port 618 nsew power bidirectional
rlabel metal4 s 296048 2128 296368 295440 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 295440 6 vssd1
port 620 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 295440 6 vssd1
port 621 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 295440 6 vssd1
port 622 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 295440 6 vssd1
port 623 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 295440 6 vssd1
port 624 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 295440 6 vssd1
port 625 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 295440 6 vssd1
port 626 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 295440 6 vssd1
port 627 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 295440 6 vssd1
port 628 nsew ground bidirectional
rlabel metal4 s 281348 2176 281668 295392 6 vccd2
port 629 nsew power bidirectional
rlabel metal4 s 250628 2176 250948 295392 6 vccd2
port 630 nsew power bidirectional
rlabel metal4 s 219908 2176 220228 295392 6 vccd2
port 631 nsew power bidirectional
rlabel metal4 s 189188 2176 189508 295392 6 vccd2
port 632 nsew power bidirectional
rlabel metal4 s 158468 2176 158788 295392 6 vccd2
port 633 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 295392 6 vccd2
port 634 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 295392 6 vccd2
port 635 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 295392 6 vccd2
port 636 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 295392 6 vccd2
port 637 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 295392 6 vccd2
port 638 nsew power bidirectional
rlabel metal4 s 265988 2176 266308 295392 6 vssd2
port 639 nsew ground bidirectional
rlabel metal4 s 235268 2176 235588 295392 6 vssd2
port 640 nsew ground bidirectional
rlabel metal4 s 204548 2176 204868 295392 6 vssd2
port 641 nsew ground bidirectional
rlabel metal4 s 173828 2176 174148 295392 6 vssd2
port 642 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 295392 6 vssd2
port 643 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 295392 6 vssd2
port 644 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 295392 6 vssd2
port 645 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 295392 6 vssd2
port 646 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 295392 6 vssd2
port 647 nsew ground bidirectional
rlabel metal4 s 282008 2176 282328 295392 6 vdda1
port 648 nsew power bidirectional
rlabel metal4 s 251288 2176 251608 295392 6 vdda1
port 649 nsew power bidirectional
rlabel metal4 s 220568 2176 220888 295392 6 vdda1
port 650 nsew power bidirectional
rlabel metal4 s 189848 2176 190168 295392 6 vdda1
port 651 nsew power bidirectional
rlabel metal4 s 159128 2176 159448 295392 6 vdda1
port 652 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 295392 6 vdda1
port 653 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 295392 6 vdda1
port 654 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 295392 6 vdda1
port 655 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 295392 6 vdda1
port 656 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 295392 6 vdda1
port 657 nsew power bidirectional
rlabel metal4 s 266648 2176 266968 295392 6 vssa1
port 658 nsew ground bidirectional
rlabel metal4 s 235928 2176 236248 295392 6 vssa1
port 659 nsew ground bidirectional
rlabel metal4 s 205208 2176 205528 295392 6 vssa1
port 660 nsew ground bidirectional
rlabel metal4 s 174488 2176 174808 295392 6 vssa1
port 661 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 295392 6 vssa1
port 662 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 295392 6 vssa1
port 663 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 295392 6 vssa1
port 664 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 295392 6 vssa1
port 665 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 295392 6 vssa1
port 666 nsew ground bidirectional
rlabel metal4 s 282668 2176 282988 295392 6 vdda2
port 667 nsew power bidirectional
rlabel metal4 s 251948 2176 252268 295392 6 vdda2
port 668 nsew power bidirectional
rlabel metal4 s 221228 2176 221548 295392 6 vdda2
port 669 nsew power bidirectional
rlabel metal4 s 190508 2176 190828 295392 6 vdda2
port 670 nsew power bidirectional
rlabel metal4 s 159788 2176 160108 295392 6 vdda2
port 671 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 295392 6 vdda2
port 672 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 295392 6 vdda2
port 673 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 295392 6 vdda2
port 674 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 295392 6 vdda2
port 675 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 295392 6 vdda2
port 676 nsew power bidirectional
rlabel metal4 s 267308 2176 267628 295392 6 vssa2
port 677 nsew ground bidirectional
rlabel metal4 s 236588 2176 236908 295392 6 vssa2
port 678 nsew ground bidirectional
rlabel metal4 s 205868 2176 206188 295392 6 vssa2
port 679 nsew ground bidirectional
rlabel metal4 s 175148 2176 175468 295392 6 vssa2
port 680 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 295392 6 vssa2
port 681 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 295392 6 vssa2
port 682 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 295392 6 vssa2
port 683 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 295392 6 vssa2
port 684 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 295392 6 vssa2
port 685 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 298000 298000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 267694638
string GDS_START 835930
<< end >>

