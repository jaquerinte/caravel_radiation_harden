VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj
  CLASS BLOCK ;
  FOREIGN user_proj ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 596.000 4.050 600.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 596.000 238.650 600.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 596.000 262.110 600.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 596.000 285.570 600.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 596.000 309.030 600.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 596.000 332.490 600.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 596.000 355.950 600.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 596.000 379.410 600.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 596.000 402.870 600.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 596.000 426.330 600.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 596.000 449.790 600.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 596.000 27.510 600.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 596.000 473.710 600.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 596.000 497.170 600.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 596.000 520.630 600.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 596.000 544.090 600.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 596.000 567.550 600.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 596.000 591.010 600.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 596.000 614.470 600.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 596.000 637.930 600.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 596.000 661.390 600.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.570 596.000 684.850 600.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 596.000 50.970 600.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 596.000 708.310 600.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 596.000 731.770 600.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.950 596.000 755.230 600.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.410 596.000 778.690 600.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 596.000 802.150 600.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.330 596.000 825.610 600.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 596.000 849.070 600.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 596.000 872.530 600.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 596.000 74.430 600.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 596.000 97.890 600.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 596.000 121.350 600.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 596.000 144.810 600.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 596.000 168.270 600.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 596.000 191.730 600.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 596.000 215.190 600.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 596.000 11.870 600.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 596.000 246.470 600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 596.000 269.930 600.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 596.000 293.390 600.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 596.000 316.850 600.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 596.000 340.310 600.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 596.000 363.770 600.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 596.000 387.230 600.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 596.000 410.690 600.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 596.000 434.150 600.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 596.000 458.070 600.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 596.000 35.330 600.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 596.000 481.530 600.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 596.000 504.990 600.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 596.000 528.450 600.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 596.000 551.910 600.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 596.000 575.370 600.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 596.000 598.830 600.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 596.000 622.290 600.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.470 596.000 645.750 600.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 596.000 669.210 600.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 596.000 692.670 600.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 596.000 58.790 600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 596.000 716.130 600.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 596.000 739.590 600.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.770 596.000 763.050 600.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.230 596.000 786.510 600.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 596.000 809.970 600.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 596.000 833.430 600.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 596.000 856.890 600.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.070 596.000 880.350 600.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 596.000 82.250 600.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 596.000 105.710 600.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 596.000 129.170 600.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 596.000 152.630 600.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 596.000 176.090 600.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 596.000 199.550 600.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 596.000 223.010 600.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 596.000 19.690 600.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 596.000 254.290 600.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 596.000 277.750 600.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 596.000 301.210 600.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 596.000 324.670 600.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 596.000 348.130 600.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 596.000 371.590 600.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 596.000 395.050 600.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 596.000 418.510 600.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 596.000 441.970 600.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 596.000 465.890 600.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 596.000 43.150 600.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 596.000 489.350 600.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.530 596.000 512.810 600.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.990 596.000 536.270 600.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 596.000 559.730 600.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 596.000 583.190 600.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 596.000 606.650 600.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 596.000 630.110 600.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 596.000 653.570 600.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 596.000 677.030 600.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 596.000 700.490 600.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 596.000 66.610 600.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.670 596.000 723.950 600.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 596.000 747.410 600.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.590 596.000 770.870 600.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 596.000 794.330 600.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.510 596.000 817.790 600.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.970 596.000 841.250 600.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.430 596.000 864.710 600.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.890 596.000 888.170 600.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 596.000 90.070 600.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 596.000 113.530 600.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 596.000 136.990 600.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 596.000 160.450 600.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 596.000 183.910 600.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 596.000 207.370 600.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 596.000 230.830 600.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 4.000 300.520 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.710 596.000 895.990 600.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 299.920 900.000 300.520 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 0.000 746.490 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.730 0.000 752.010 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.250 0.000 757.530 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.770 0.000 763.050 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.290 0.000 768.570 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.810 0.000 774.090 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 0.000 785.130 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.370 0.000 790.650 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 0.000 796.170 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.410 0.000 801.690 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.930 0.000 807.210 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.450 0.000 812.730 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.490 0.000 823.770 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 0.000 829.290 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.530 0.000 834.810 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.050 0.000 840.330 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.570 0.000 845.850 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.090 0.000 851.370 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 0.000 856.890 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.130 0.000 862.410 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.650 0.000 867.930 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.170 0.000 873.450 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.690 0.000 878.970 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.210 0.000 884.490 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.730 0.000 890.010 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 0.000 895.530 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 0.000 305.350 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 0.000 349.510 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 0.000 360.550 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 0.000 366.070 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 0.000 382.630 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 0.000 399.190 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 0.000 410.230 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 0.000 421.270 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 0.000 432.310 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 0.000 448.870 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 0.000 459.910 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.150 0.000 465.430 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 0.000 470.950 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 0.000 476.470 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 0.000 487.510 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.270 0.000 498.550 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 0.000 520.630 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 0.000 526.150 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 0.000 548.230 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 0.000 553.750 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 0.000 559.270 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 0.000 564.790 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 0.000 575.830 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 0.000 581.350 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 0.000 586.870 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 0.000 592.390 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 0.000 597.910 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 0.000 602.970 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.210 0.000 608.490 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.730 0.000 614.010 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.250 0.000 619.530 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 0.000 630.570 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.810 0.000 636.090 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 0.000 641.610 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.850 0.000 647.130 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 0.000 652.650 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 0.000 658.170 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 0.000 669.210 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 0.000 674.730 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 0.000 680.250 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 0.000 685.770 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.010 0.000 691.290 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.530 0.000 696.810 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 0.000 702.330 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 0.000 707.850 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 0.000 713.370 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 0.000 718.890 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 0.000 724.410 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 0.000 735.450 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 0.000 748.330 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 0.000 759.370 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.610 0.000 764.890 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.130 0.000 770.410 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 0.000 775.930 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 0.000 781.450 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 0.000 786.970 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 0.000 798.010 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.250 0.000 803.530 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.770 0.000 809.050 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 0.000 814.570 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 0.000 820.090 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.330 0.000 825.610 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.370 0.000 836.650 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 0.000 842.170 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.410 0.000 847.690 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.930 0.000 853.210 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.450 0.000 858.730 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.970 0.000 864.250 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 0.000 869.770 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 0.000 875.290 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.530 0.000 880.810 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.050 0.000 886.330 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.570 0.000 891.850 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.090 0.000 897.370 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 0.000 334.790 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 0.000 384.470 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 0.000 395.510 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 0.000 401.030 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 0.000 412.070 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 0.000 423.110 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 0.000 434.150 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.910 0.000 445.190 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 0.000 450.710 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 0.000 456.230 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 0.000 472.790 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 0.000 478.310 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 0.000 483.830 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 0.000 494.870 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.110 0.000 500.390 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 0.000 511.430 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 0.000 516.950 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 0.000 527.990 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 0.000 533.510 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 0.000 539.030 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 0.000 550.070 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 0.000 555.590 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 0.000 561.110 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 0.000 566.630 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 0.000 572.150 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 0.000 577.670 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 0.000 588.710 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 0.000 594.230 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 0.000 604.810 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.050 0.000 610.330 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 0.000 621.370 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 0.000 626.890 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 0.000 632.410 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 0.000 643.450 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 0.000 648.970 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 0.000 654.490 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 0.000 660.010 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 0.000 665.530 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 0.000 671.050 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 0.000 682.090 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 0.000 687.610 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 0.000 693.130 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.370 0.000 698.650 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 0.000 704.170 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 0.000 709.690 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 0.000 720.730 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.970 0.000 726.250 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 0.000 731.770 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 0.000 737.290 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 0.000 742.810 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.410 0.000 755.690 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.930 0.000 761.210 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 0.000 772.250 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.490 0.000 777.770 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 0.000 783.290 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.530 0.000 788.810 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 0.000 794.330 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.570 0.000 799.850 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 0.000 805.370 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.610 0.000 810.890 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.130 0.000 816.410 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.650 0.000 821.930 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.170 0.000 827.450 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.690 0.000 832.970 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.210 0.000 838.490 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 0.000 844.010 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.250 0.000 849.530 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.770 0.000 855.050 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 0.000 860.570 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.810 0.000 866.090 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.330 0.000 871.610 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.850 0.000 877.130 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 0.000 882.650 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.890 0.000 888.170 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.410 0.000 893.690 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.930 0.000 899.210 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 0.000 303.510 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 0.000 353.190 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 0.000 435.990 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 0.000 463.590 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.830 0.000 469.110 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 0.000 513.270 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 0.000 524.310 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 0.000 535.350 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 0.000 540.870 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 0.000 551.910 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 0.000 568.470 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 0.000 573.990 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 0.000 579.510 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 0.000 585.030 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.270 0.000 590.550 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 0.000 601.130 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 0.000 606.650 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 0.000 617.690 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 0.000 623.210 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.970 0.000 634.250 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 0.000 639.770 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 0.000 645.290 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 0.000 656.330 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.570 0.000 661.850 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 0.000 672.890 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.130 0.000 678.410 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.650 0.000 683.930 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.690 0.000 694.970 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.730 0.000 706.010 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 0.000 711.530 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 0.000 717.050 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 0.000 722.570 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 0.000 733.610 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.850 0.000 739.130 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.370 0.000 744.650 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END la_oenb[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 0.000 0.830 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 792.340 10.880 793.940 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 587.520 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 869.140 10.880 870.740 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 715.540 10.880 717.140 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 587.520 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 795.640 10.880 797.240 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 642.040 10.880 643.640 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.440 10.880 490.040 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 587.520 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 872.440 10.880 874.040 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 718.840 10.880 720.440 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 565.240 10.880 566.840 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.640 10.880 413.240 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 587.520 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 798.940 10.880 800.540 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 645.340 10.880 646.940 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.740 10.880 493.340 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 587.520 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 875.740 10.880 877.340 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 722.140 10.880 723.740 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.540 10.880 570.140 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.940 10.880 416.540 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 587.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 0.530 6.840 899.230 587.760 ;
      LAYER met2 ;
        RECT 0.560 595.720 3.490 596.000 ;
        RECT 4.330 595.720 11.310 596.000 ;
        RECT 12.150 595.720 19.130 596.000 ;
        RECT 19.970 595.720 26.950 596.000 ;
        RECT 27.790 595.720 34.770 596.000 ;
        RECT 35.610 595.720 42.590 596.000 ;
        RECT 43.430 595.720 50.410 596.000 ;
        RECT 51.250 595.720 58.230 596.000 ;
        RECT 59.070 595.720 66.050 596.000 ;
        RECT 66.890 595.720 73.870 596.000 ;
        RECT 74.710 595.720 81.690 596.000 ;
        RECT 82.530 595.720 89.510 596.000 ;
        RECT 90.350 595.720 97.330 596.000 ;
        RECT 98.170 595.720 105.150 596.000 ;
        RECT 105.990 595.720 112.970 596.000 ;
        RECT 113.810 595.720 120.790 596.000 ;
        RECT 121.630 595.720 128.610 596.000 ;
        RECT 129.450 595.720 136.430 596.000 ;
        RECT 137.270 595.720 144.250 596.000 ;
        RECT 145.090 595.720 152.070 596.000 ;
        RECT 152.910 595.720 159.890 596.000 ;
        RECT 160.730 595.720 167.710 596.000 ;
        RECT 168.550 595.720 175.530 596.000 ;
        RECT 176.370 595.720 183.350 596.000 ;
        RECT 184.190 595.720 191.170 596.000 ;
        RECT 192.010 595.720 198.990 596.000 ;
        RECT 199.830 595.720 206.810 596.000 ;
        RECT 207.650 595.720 214.630 596.000 ;
        RECT 215.470 595.720 222.450 596.000 ;
        RECT 223.290 595.720 230.270 596.000 ;
        RECT 231.110 595.720 238.090 596.000 ;
        RECT 238.930 595.720 245.910 596.000 ;
        RECT 246.750 595.720 253.730 596.000 ;
        RECT 254.570 595.720 261.550 596.000 ;
        RECT 262.390 595.720 269.370 596.000 ;
        RECT 270.210 595.720 277.190 596.000 ;
        RECT 278.030 595.720 285.010 596.000 ;
        RECT 285.850 595.720 292.830 596.000 ;
        RECT 293.670 595.720 300.650 596.000 ;
        RECT 301.490 595.720 308.470 596.000 ;
        RECT 309.310 595.720 316.290 596.000 ;
        RECT 317.130 595.720 324.110 596.000 ;
        RECT 324.950 595.720 331.930 596.000 ;
        RECT 332.770 595.720 339.750 596.000 ;
        RECT 340.590 595.720 347.570 596.000 ;
        RECT 348.410 595.720 355.390 596.000 ;
        RECT 356.230 595.720 363.210 596.000 ;
        RECT 364.050 595.720 371.030 596.000 ;
        RECT 371.870 595.720 378.850 596.000 ;
        RECT 379.690 595.720 386.670 596.000 ;
        RECT 387.510 595.720 394.490 596.000 ;
        RECT 395.330 595.720 402.310 596.000 ;
        RECT 403.150 595.720 410.130 596.000 ;
        RECT 410.970 595.720 417.950 596.000 ;
        RECT 418.790 595.720 425.770 596.000 ;
        RECT 426.610 595.720 433.590 596.000 ;
        RECT 434.430 595.720 441.410 596.000 ;
        RECT 442.250 595.720 449.230 596.000 ;
        RECT 450.070 595.720 457.510 596.000 ;
        RECT 458.350 595.720 465.330 596.000 ;
        RECT 466.170 595.720 473.150 596.000 ;
        RECT 473.990 595.720 480.970 596.000 ;
        RECT 481.810 595.720 488.790 596.000 ;
        RECT 489.630 595.720 496.610 596.000 ;
        RECT 497.450 595.720 504.430 596.000 ;
        RECT 505.270 595.720 512.250 596.000 ;
        RECT 513.090 595.720 520.070 596.000 ;
        RECT 520.910 595.720 527.890 596.000 ;
        RECT 528.730 595.720 535.710 596.000 ;
        RECT 536.550 595.720 543.530 596.000 ;
        RECT 544.370 595.720 551.350 596.000 ;
        RECT 552.190 595.720 559.170 596.000 ;
        RECT 560.010 595.720 566.990 596.000 ;
        RECT 567.830 595.720 574.810 596.000 ;
        RECT 575.650 595.720 582.630 596.000 ;
        RECT 583.470 595.720 590.450 596.000 ;
        RECT 591.290 595.720 598.270 596.000 ;
        RECT 599.110 595.720 606.090 596.000 ;
        RECT 606.930 595.720 613.910 596.000 ;
        RECT 614.750 595.720 621.730 596.000 ;
        RECT 622.570 595.720 629.550 596.000 ;
        RECT 630.390 595.720 637.370 596.000 ;
        RECT 638.210 595.720 645.190 596.000 ;
        RECT 646.030 595.720 653.010 596.000 ;
        RECT 653.850 595.720 660.830 596.000 ;
        RECT 661.670 595.720 668.650 596.000 ;
        RECT 669.490 595.720 676.470 596.000 ;
        RECT 677.310 595.720 684.290 596.000 ;
        RECT 685.130 595.720 692.110 596.000 ;
        RECT 692.950 595.720 699.930 596.000 ;
        RECT 700.770 595.720 707.750 596.000 ;
        RECT 708.590 595.720 715.570 596.000 ;
        RECT 716.410 595.720 723.390 596.000 ;
        RECT 724.230 595.720 731.210 596.000 ;
        RECT 732.050 595.720 739.030 596.000 ;
        RECT 739.870 595.720 746.850 596.000 ;
        RECT 747.690 595.720 754.670 596.000 ;
        RECT 755.510 595.720 762.490 596.000 ;
        RECT 763.330 595.720 770.310 596.000 ;
        RECT 771.150 595.720 778.130 596.000 ;
        RECT 778.970 595.720 785.950 596.000 ;
        RECT 786.790 595.720 793.770 596.000 ;
        RECT 794.610 595.720 801.590 596.000 ;
        RECT 802.430 595.720 809.410 596.000 ;
        RECT 810.250 595.720 817.230 596.000 ;
        RECT 818.070 595.720 825.050 596.000 ;
        RECT 825.890 595.720 832.870 596.000 ;
        RECT 833.710 595.720 840.690 596.000 ;
        RECT 841.530 595.720 848.510 596.000 ;
        RECT 849.350 595.720 856.330 596.000 ;
        RECT 857.170 595.720 864.150 596.000 ;
        RECT 864.990 595.720 871.970 596.000 ;
        RECT 872.810 595.720 879.790 596.000 ;
        RECT 880.630 595.720 887.610 596.000 ;
        RECT 888.450 595.720 895.430 596.000 ;
        RECT 896.270 595.720 899.200 596.000 ;
        RECT 0.560 4.280 899.200 595.720 ;
        RECT 1.110 4.000 1.650 4.280 ;
        RECT 2.490 4.000 3.490 4.280 ;
        RECT 4.330 4.000 5.330 4.280 ;
        RECT 6.170 4.000 7.170 4.280 ;
        RECT 8.010 4.000 9.010 4.280 ;
        RECT 9.850 4.000 10.850 4.280 ;
        RECT 11.690 4.000 12.690 4.280 ;
        RECT 13.530 4.000 14.530 4.280 ;
        RECT 15.370 4.000 16.370 4.280 ;
        RECT 17.210 4.000 18.210 4.280 ;
        RECT 19.050 4.000 20.050 4.280 ;
        RECT 20.890 4.000 21.890 4.280 ;
        RECT 22.730 4.000 23.730 4.280 ;
        RECT 24.570 4.000 25.570 4.280 ;
        RECT 26.410 4.000 27.410 4.280 ;
        RECT 28.250 4.000 29.250 4.280 ;
        RECT 30.090 4.000 31.090 4.280 ;
        RECT 31.930 4.000 32.930 4.280 ;
        RECT 33.770 4.000 34.770 4.280 ;
        RECT 35.610 4.000 36.610 4.280 ;
        RECT 37.450 4.000 38.450 4.280 ;
        RECT 39.290 4.000 40.290 4.280 ;
        RECT 41.130 4.000 42.130 4.280 ;
        RECT 42.970 4.000 43.970 4.280 ;
        RECT 44.810 4.000 45.810 4.280 ;
        RECT 46.650 4.000 47.650 4.280 ;
        RECT 48.490 4.000 49.490 4.280 ;
        RECT 50.330 4.000 51.330 4.280 ;
        RECT 52.170 4.000 53.170 4.280 ;
        RECT 54.010 4.000 55.010 4.280 ;
        RECT 55.850 4.000 56.850 4.280 ;
        RECT 57.690 4.000 58.690 4.280 ;
        RECT 59.530 4.000 60.530 4.280 ;
        RECT 61.370 4.000 62.370 4.280 ;
        RECT 63.210 4.000 64.210 4.280 ;
        RECT 65.050 4.000 66.050 4.280 ;
        RECT 66.890 4.000 67.890 4.280 ;
        RECT 68.730 4.000 69.730 4.280 ;
        RECT 70.570 4.000 71.570 4.280 ;
        RECT 72.410 4.000 73.410 4.280 ;
        RECT 74.250 4.000 75.250 4.280 ;
        RECT 76.090 4.000 77.090 4.280 ;
        RECT 77.930 4.000 78.930 4.280 ;
        RECT 79.770 4.000 80.770 4.280 ;
        RECT 81.610 4.000 82.610 4.280 ;
        RECT 83.450 4.000 84.450 4.280 ;
        RECT 85.290 4.000 86.290 4.280 ;
        RECT 87.130 4.000 88.130 4.280 ;
        RECT 88.970 4.000 89.970 4.280 ;
        RECT 90.810 4.000 91.810 4.280 ;
        RECT 92.650 4.000 93.650 4.280 ;
        RECT 94.490 4.000 95.490 4.280 ;
        RECT 96.330 4.000 97.330 4.280 ;
        RECT 98.170 4.000 99.170 4.280 ;
        RECT 100.010 4.000 101.010 4.280 ;
        RECT 101.850 4.000 102.850 4.280 ;
        RECT 103.690 4.000 104.690 4.280 ;
        RECT 105.530 4.000 106.530 4.280 ;
        RECT 107.370 4.000 108.370 4.280 ;
        RECT 109.210 4.000 110.210 4.280 ;
        RECT 111.050 4.000 112.050 4.280 ;
        RECT 112.890 4.000 113.890 4.280 ;
        RECT 114.730 4.000 115.730 4.280 ;
        RECT 116.570 4.000 117.570 4.280 ;
        RECT 118.410 4.000 119.410 4.280 ;
        RECT 120.250 4.000 121.250 4.280 ;
        RECT 122.090 4.000 123.090 4.280 ;
        RECT 123.930 4.000 124.930 4.280 ;
        RECT 125.770 4.000 126.770 4.280 ;
        RECT 127.610 4.000 128.610 4.280 ;
        RECT 129.450 4.000 130.450 4.280 ;
        RECT 131.290 4.000 132.290 4.280 ;
        RECT 133.130 4.000 134.130 4.280 ;
        RECT 134.970 4.000 135.970 4.280 ;
        RECT 136.810 4.000 137.810 4.280 ;
        RECT 138.650 4.000 139.650 4.280 ;
        RECT 140.490 4.000 141.490 4.280 ;
        RECT 142.330 4.000 143.330 4.280 ;
        RECT 144.170 4.000 145.170 4.280 ;
        RECT 146.010 4.000 147.010 4.280 ;
        RECT 147.850 4.000 148.850 4.280 ;
        RECT 149.690 4.000 150.690 4.280 ;
        RECT 151.530 4.000 152.530 4.280 ;
        RECT 153.370 4.000 154.370 4.280 ;
        RECT 155.210 4.000 156.210 4.280 ;
        RECT 157.050 4.000 158.050 4.280 ;
        RECT 158.890 4.000 159.890 4.280 ;
        RECT 160.730 4.000 161.730 4.280 ;
        RECT 162.570 4.000 163.570 4.280 ;
        RECT 164.410 4.000 165.410 4.280 ;
        RECT 166.250 4.000 167.250 4.280 ;
        RECT 168.090 4.000 169.090 4.280 ;
        RECT 169.930 4.000 170.930 4.280 ;
        RECT 171.770 4.000 172.770 4.280 ;
        RECT 173.610 4.000 174.610 4.280 ;
        RECT 175.450 4.000 176.450 4.280 ;
        RECT 177.290 4.000 178.290 4.280 ;
        RECT 179.130 4.000 180.130 4.280 ;
        RECT 180.970 4.000 181.970 4.280 ;
        RECT 182.810 4.000 183.810 4.280 ;
        RECT 184.650 4.000 185.650 4.280 ;
        RECT 186.490 4.000 187.490 4.280 ;
        RECT 188.330 4.000 189.330 4.280 ;
        RECT 190.170 4.000 191.170 4.280 ;
        RECT 192.010 4.000 193.010 4.280 ;
        RECT 193.850 4.000 194.850 4.280 ;
        RECT 195.690 4.000 196.690 4.280 ;
        RECT 197.530 4.000 198.530 4.280 ;
        RECT 199.370 4.000 200.370 4.280 ;
        RECT 201.210 4.000 202.210 4.280 ;
        RECT 203.050 4.000 204.050 4.280 ;
        RECT 204.890 4.000 205.890 4.280 ;
        RECT 206.730 4.000 207.730 4.280 ;
        RECT 208.570 4.000 209.570 4.280 ;
        RECT 210.410 4.000 211.410 4.280 ;
        RECT 212.250 4.000 213.250 4.280 ;
        RECT 214.090 4.000 215.090 4.280 ;
        RECT 215.930 4.000 216.930 4.280 ;
        RECT 217.770 4.000 218.770 4.280 ;
        RECT 219.610 4.000 220.610 4.280 ;
        RECT 221.450 4.000 222.450 4.280 ;
        RECT 223.290 4.000 224.290 4.280 ;
        RECT 225.130 4.000 226.130 4.280 ;
        RECT 226.970 4.000 227.970 4.280 ;
        RECT 228.810 4.000 229.810 4.280 ;
        RECT 230.650 4.000 231.650 4.280 ;
        RECT 232.490 4.000 233.490 4.280 ;
        RECT 234.330 4.000 235.330 4.280 ;
        RECT 236.170 4.000 237.170 4.280 ;
        RECT 238.010 4.000 239.010 4.280 ;
        RECT 239.850 4.000 240.850 4.280 ;
        RECT 241.690 4.000 242.690 4.280 ;
        RECT 243.530 4.000 244.530 4.280 ;
        RECT 245.370 4.000 246.370 4.280 ;
        RECT 247.210 4.000 248.210 4.280 ;
        RECT 249.050 4.000 250.050 4.280 ;
        RECT 250.890 4.000 251.890 4.280 ;
        RECT 252.730 4.000 253.730 4.280 ;
        RECT 254.570 4.000 255.570 4.280 ;
        RECT 256.410 4.000 257.410 4.280 ;
        RECT 258.250 4.000 259.250 4.280 ;
        RECT 260.090 4.000 261.090 4.280 ;
        RECT 261.930 4.000 262.930 4.280 ;
        RECT 263.770 4.000 264.770 4.280 ;
        RECT 265.610 4.000 266.610 4.280 ;
        RECT 267.450 4.000 268.450 4.280 ;
        RECT 269.290 4.000 270.290 4.280 ;
        RECT 271.130 4.000 272.130 4.280 ;
        RECT 272.970 4.000 273.970 4.280 ;
        RECT 274.810 4.000 275.810 4.280 ;
        RECT 276.650 4.000 277.650 4.280 ;
        RECT 278.490 4.000 279.490 4.280 ;
        RECT 280.330 4.000 281.330 4.280 ;
        RECT 282.170 4.000 283.170 4.280 ;
        RECT 284.010 4.000 285.010 4.280 ;
        RECT 285.850 4.000 286.850 4.280 ;
        RECT 287.690 4.000 288.690 4.280 ;
        RECT 289.530 4.000 290.530 4.280 ;
        RECT 291.370 4.000 292.370 4.280 ;
        RECT 293.210 4.000 294.210 4.280 ;
        RECT 295.050 4.000 296.050 4.280 ;
        RECT 296.890 4.000 297.890 4.280 ;
        RECT 298.730 4.000 299.730 4.280 ;
        RECT 300.570 4.000 301.110 4.280 ;
        RECT 301.950 4.000 302.950 4.280 ;
        RECT 303.790 4.000 304.790 4.280 ;
        RECT 305.630 4.000 306.630 4.280 ;
        RECT 307.470 4.000 308.470 4.280 ;
        RECT 309.310 4.000 310.310 4.280 ;
        RECT 311.150 4.000 312.150 4.280 ;
        RECT 312.990 4.000 313.990 4.280 ;
        RECT 314.830 4.000 315.830 4.280 ;
        RECT 316.670 4.000 317.670 4.280 ;
        RECT 318.510 4.000 319.510 4.280 ;
        RECT 320.350 4.000 321.350 4.280 ;
        RECT 322.190 4.000 323.190 4.280 ;
        RECT 324.030 4.000 325.030 4.280 ;
        RECT 325.870 4.000 326.870 4.280 ;
        RECT 327.710 4.000 328.710 4.280 ;
        RECT 329.550 4.000 330.550 4.280 ;
        RECT 331.390 4.000 332.390 4.280 ;
        RECT 333.230 4.000 334.230 4.280 ;
        RECT 335.070 4.000 336.070 4.280 ;
        RECT 336.910 4.000 337.910 4.280 ;
        RECT 338.750 4.000 339.750 4.280 ;
        RECT 340.590 4.000 341.590 4.280 ;
        RECT 342.430 4.000 343.430 4.280 ;
        RECT 344.270 4.000 345.270 4.280 ;
        RECT 346.110 4.000 347.110 4.280 ;
        RECT 347.950 4.000 348.950 4.280 ;
        RECT 349.790 4.000 350.790 4.280 ;
        RECT 351.630 4.000 352.630 4.280 ;
        RECT 353.470 4.000 354.470 4.280 ;
        RECT 355.310 4.000 356.310 4.280 ;
        RECT 357.150 4.000 358.150 4.280 ;
        RECT 358.990 4.000 359.990 4.280 ;
        RECT 360.830 4.000 361.830 4.280 ;
        RECT 362.670 4.000 363.670 4.280 ;
        RECT 364.510 4.000 365.510 4.280 ;
        RECT 366.350 4.000 367.350 4.280 ;
        RECT 368.190 4.000 369.190 4.280 ;
        RECT 370.030 4.000 371.030 4.280 ;
        RECT 371.870 4.000 372.870 4.280 ;
        RECT 373.710 4.000 374.710 4.280 ;
        RECT 375.550 4.000 376.550 4.280 ;
        RECT 377.390 4.000 378.390 4.280 ;
        RECT 379.230 4.000 380.230 4.280 ;
        RECT 381.070 4.000 382.070 4.280 ;
        RECT 382.910 4.000 383.910 4.280 ;
        RECT 384.750 4.000 385.750 4.280 ;
        RECT 386.590 4.000 387.590 4.280 ;
        RECT 388.430 4.000 389.430 4.280 ;
        RECT 390.270 4.000 391.270 4.280 ;
        RECT 392.110 4.000 393.110 4.280 ;
        RECT 393.950 4.000 394.950 4.280 ;
        RECT 395.790 4.000 396.790 4.280 ;
        RECT 397.630 4.000 398.630 4.280 ;
        RECT 399.470 4.000 400.470 4.280 ;
        RECT 401.310 4.000 402.310 4.280 ;
        RECT 403.150 4.000 404.150 4.280 ;
        RECT 404.990 4.000 405.990 4.280 ;
        RECT 406.830 4.000 407.830 4.280 ;
        RECT 408.670 4.000 409.670 4.280 ;
        RECT 410.510 4.000 411.510 4.280 ;
        RECT 412.350 4.000 413.350 4.280 ;
        RECT 414.190 4.000 415.190 4.280 ;
        RECT 416.030 4.000 417.030 4.280 ;
        RECT 417.870 4.000 418.870 4.280 ;
        RECT 419.710 4.000 420.710 4.280 ;
        RECT 421.550 4.000 422.550 4.280 ;
        RECT 423.390 4.000 424.390 4.280 ;
        RECT 425.230 4.000 426.230 4.280 ;
        RECT 427.070 4.000 428.070 4.280 ;
        RECT 428.910 4.000 429.910 4.280 ;
        RECT 430.750 4.000 431.750 4.280 ;
        RECT 432.590 4.000 433.590 4.280 ;
        RECT 434.430 4.000 435.430 4.280 ;
        RECT 436.270 4.000 437.270 4.280 ;
        RECT 438.110 4.000 439.110 4.280 ;
        RECT 439.950 4.000 440.950 4.280 ;
        RECT 441.790 4.000 442.790 4.280 ;
        RECT 443.630 4.000 444.630 4.280 ;
        RECT 445.470 4.000 446.470 4.280 ;
        RECT 447.310 4.000 448.310 4.280 ;
        RECT 449.150 4.000 450.150 4.280 ;
        RECT 450.990 4.000 451.990 4.280 ;
        RECT 452.830 4.000 453.830 4.280 ;
        RECT 454.670 4.000 455.670 4.280 ;
        RECT 456.510 4.000 457.510 4.280 ;
        RECT 458.350 4.000 459.350 4.280 ;
        RECT 460.190 4.000 461.190 4.280 ;
        RECT 462.030 4.000 463.030 4.280 ;
        RECT 463.870 4.000 464.870 4.280 ;
        RECT 465.710 4.000 466.710 4.280 ;
        RECT 467.550 4.000 468.550 4.280 ;
        RECT 469.390 4.000 470.390 4.280 ;
        RECT 471.230 4.000 472.230 4.280 ;
        RECT 473.070 4.000 474.070 4.280 ;
        RECT 474.910 4.000 475.910 4.280 ;
        RECT 476.750 4.000 477.750 4.280 ;
        RECT 478.590 4.000 479.590 4.280 ;
        RECT 480.430 4.000 481.430 4.280 ;
        RECT 482.270 4.000 483.270 4.280 ;
        RECT 484.110 4.000 485.110 4.280 ;
        RECT 485.950 4.000 486.950 4.280 ;
        RECT 487.790 4.000 488.790 4.280 ;
        RECT 489.630 4.000 490.630 4.280 ;
        RECT 491.470 4.000 492.470 4.280 ;
        RECT 493.310 4.000 494.310 4.280 ;
        RECT 495.150 4.000 496.150 4.280 ;
        RECT 496.990 4.000 497.990 4.280 ;
        RECT 498.830 4.000 499.830 4.280 ;
        RECT 500.670 4.000 501.670 4.280 ;
        RECT 502.510 4.000 503.510 4.280 ;
        RECT 504.350 4.000 505.350 4.280 ;
        RECT 506.190 4.000 507.190 4.280 ;
        RECT 508.030 4.000 509.030 4.280 ;
        RECT 509.870 4.000 510.870 4.280 ;
        RECT 511.710 4.000 512.710 4.280 ;
        RECT 513.550 4.000 514.550 4.280 ;
        RECT 515.390 4.000 516.390 4.280 ;
        RECT 517.230 4.000 518.230 4.280 ;
        RECT 519.070 4.000 520.070 4.280 ;
        RECT 520.910 4.000 521.910 4.280 ;
        RECT 522.750 4.000 523.750 4.280 ;
        RECT 524.590 4.000 525.590 4.280 ;
        RECT 526.430 4.000 527.430 4.280 ;
        RECT 528.270 4.000 529.270 4.280 ;
        RECT 530.110 4.000 531.110 4.280 ;
        RECT 531.950 4.000 532.950 4.280 ;
        RECT 533.790 4.000 534.790 4.280 ;
        RECT 535.630 4.000 536.630 4.280 ;
        RECT 537.470 4.000 538.470 4.280 ;
        RECT 539.310 4.000 540.310 4.280 ;
        RECT 541.150 4.000 542.150 4.280 ;
        RECT 542.990 4.000 543.990 4.280 ;
        RECT 544.830 4.000 545.830 4.280 ;
        RECT 546.670 4.000 547.670 4.280 ;
        RECT 548.510 4.000 549.510 4.280 ;
        RECT 550.350 4.000 551.350 4.280 ;
        RECT 552.190 4.000 553.190 4.280 ;
        RECT 554.030 4.000 555.030 4.280 ;
        RECT 555.870 4.000 556.870 4.280 ;
        RECT 557.710 4.000 558.710 4.280 ;
        RECT 559.550 4.000 560.550 4.280 ;
        RECT 561.390 4.000 562.390 4.280 ;
        RECT 563.230 4.000 564.230 4.280 ;
        RECT 565.070 4.000 566.070 4.280 ;
        RECT 566.910 4.000 567.910 4.280 ;
        RECT 568.750 4.000 569.750 4.280 ;
        RECT 570.590 4.000 571.590 4.280 ;
        RECT 572.430 4.000 573.430 4.280 ;
        RECT 574.270 4.000 575.270 4.280 ;
        RECT 576.110 4.000 577.110 4.280 ;
        RECT 577.950 4.000 578.950 4.280 ;
        RECT 579.790 4.000 580.790 4.280 ;
        RECT 581.630 4.000 582.630 4.280 ;
        RECT 583.470 4.000 584.470 4.280 ;
        RECT 585.310 4.000 586.310 4.280 ;
        RECT 587.150 4.000 588.150 4.280 ;
        RECT 588.990 4.000 589.990 4.280 ;
        RECT 590.830 4.000 591.830 4.280 ;
        RECT 592.670 4.000 593.670 4.280 ;
        RECT 594.510 4.000 595.510 4.280 ;
        RECT 596.350 4.000 597.350 4.280 ;
        RECT 598.190 4.000 599.190 4.280 ;
        RECT 600.030 4.000 600.570 4.280 ;
        RECT 601.410 4.000 602.410 4.280 ;
        RECT 603.250 4.000 604.250 4.280 ;
        RECT 605.090 4.000 606.090 4.280 ;
        RECT 606.930 4.000 607.930 4.280 ;
        RECT 608.770 4.000 609.770 4.280 ;
        RECT 610.610 4.000 611.610 4.280 ;
        RECT 612.450 4.000 613.450 4.280 ;
        RECT 614.290 4.000 615.290 4.280 ;
        RECT 616.130 4.000 617.130 4.280 ;
        RECT 617.970 4.000 618.970 4.280 ;
        RECT 619.810 4.000 620.810 4.280 ;
        RECT 621.650 4.000 622.650 4.280 ;
        RECT 623.490 4.000 624.490 4.280 ;
        RECT 625.330 4.000 626.330 4.280 ;
        RECT 627.170 4.000 628.170 4.280 ;
        RECT 629.010 4.000 630.010 4.280 ;
        RECT 630.850 4.000 631.850 4.280 ;
        RECT 632.690 4.000 633.690 4.280 ;
        RECT 634.530 4.000 635.530 4.280 ;
        RECT 636.370 4.000 637.370 4.280 ;
        RECT 638.210 4.000 639.210 4.280 ;
        RECT 640.050 4.000 641.050 4.280 ;
        RECT 641.890 4.000 642.890 4.280 ;
        RECT 643.730 4.000 644.730 4.280 ;
        RECT 645.570 4.000 646.570 4.280 ;
        RECT 647.410 4.000 648.410 4.280 ;
        RECT 649.250 4.000 650.250 4.280 ;
        RECT 651.090 4.000 652.090 4.280 ;
        RECT 652.930 4.000 653.930 4.280 ;
        RECT 654.770 4.000 655.770 4.280 ;
        RECT 656.610 4.000 657.610 4.280 ;
        RECT 658.450 4.000 659.450 4.280 ;
        RECT 660.290 4.000 661.290 4.280 ;
        RECT 662.130 4.000 663.130 4.280 ;
        RECT 663.970 4.000 664.970 4.280 ;
        RECT 665.810 4.000 666.810 4.280 ;
        RECT 667.650 4.000 668.650 4.280 ;
        RECT 669.490 4.000 670.490 4.280 ;
        RECT 671.330 4.000 672.330 4.280 ;
        RECT 673.170 4.000 674.170 4.280 ;
        RECT 675.010 4.000 676.010 4.280 ;
        RECT 676.850 4.000 677.850 4.280 ;
        RECT 678.690 4.000 679.690 4.280 ;
        RECT 680.530 4.000 681.530 4.280 ;
        RECT 682.370 4.000 683.370 4.280 ;
        RECT 684.210 4.000 685.210 4.280 ;
        RECT 686.050 4.000 687.050 4.280 ;
        RECT 687.890 4.000 688.890 4.280 ;
        RECT 689.730 4.000 690.730 4.280 ;
        RECT 691.570 4.000 692.570 4.280 ;
        RECT 693.410 4.000 694.410 4.280 ;
        RECT 695.250 4.000 696.250 4.280 ;
        RECT 697.090 4.000 698.090 4.280 ;
        RECT 698.930 4.000 699.930 4.280 ;
        RECT 700.770 4.000 701.770 4.280 ;
        RECT 702.610 4.000 703.610 4.280 ;
        RECT 704.450 4.000 705.450 4.280 ;
        RECT 706.290 4.000 707.290 4.280 ;
        RECT 708.130 4.000 709.130 4.280 ;
        RECT 709.970 4.000 710.970 4.280 ;
        RECT 711.810 4.000 712.810 4.280 ;
        RECT 713.650 4.000 714.650 4.280 ;
        RECT 715.490 4.000 716.490 4.280 ;
        RECT 717.330 4.000 718.330 4.280 ;
        RECT 719.170 4.000 720.170 4.280 ;
        RECT 721.010 4.000 722.010 4.280 ;
        RECT 722.850 4.000 723.850 4.280 ;
        RECT 724.690 4.000 725.690 4.280 ;
        RECT 726.530 4.000 727.530 4.280 ;
        RECT 728.370 4.000 729.370 4.280 ;
        RECT 730.210 4.000 731.210 4.280 ;
        RECT 732.050 4.000 733.050 4.280 ;
        RECT 733.890 4.000 734.890 4.280 ;
        RECT 735.730 4.000 736.730 4.280 ;
        RECT 737.570 4.000 738.570 4.280 ;
        RECT 739.410 4.000 740.410 4.280 ;
        RECT 741.250 4.000 742.250 4.280 ;
        RECT 743.090 4.000 744.090 4.280 ;
        RECT 744.930 4.000 745.930 4.280 ;
        RECT 746.770 4.000 747.770 4.280 ;
        RECT 748.610 4.000 749.610 4.280 ;
        RECT 750.450 4.000 751.450 4.280 ;
        RECT 752.290 4.000 753.290 4.280 ;
        RECT 754.130 4.000 755.130 4.280 ;
        RECT 755.970 4.000 756.970 4.280 ;
        RECT 757.810 4.000 758.810 4.280 ;
        RECT 759.650 4.000 760.650 4.280 ;
        RECT 761.490 4.000 762.490 4.280 ;
        RECT 763.330 4.000 764.330 4.280 ;
        RECT 765.170 4.000 766.170 4.280 ;
        RECT 767.010 4.000 768.010 4.280 ;
        RECT 768.850 4.000 769.850 4.280 ;
        RECT 770.690 4.000 771.690 4.280 ;
        RECT 772.530 4.000 773.530 4.280 ;
        RECT 774.370 4.000 775.370 4.280 ;
        RECT 776.210 4.000 777.210 4.280 ;
        RECT 778.050 4.000 779.050 4.280 ;
        RECT 779.890 4.000 780.890 4.280 ;
        RECT 781.730 4.000 782.730 4.280 ;
        RECT 783.570 4.000 784.570 4.280 ;
        RECT 785.410 4.000 786.410 4.280 ;
        RECT 787.250 4.000 788.250 4.280 ;
        RECT 789.090 4.000 790.090 4.280 ;
        RECT 790.930 4.000 791.930 4.280 ;
        RECT 792.770 4.000 793.770 4.280 ;
        RECT 794.610 4.000 795.610 4.280 ;
        RECT 796.450 4.000 797.450 4.280 ;
        RECT 798.290 4.000 799.290 4.280 ;
        RECT 800.130 4.000 801.130 4.280 ;
        RECT 801.970 4.000 802.970 4.280 ;
        RECT 803.810 4.000 804.810 4.280 ;
        RECT 805.650 4.000 806.650 4.280 ;
        RECT 807.490 4.000 808.490 4.280 ;
        RECT 809.330 4.000 810.330 4.280 ;
        RECT 811.170 4.000 812.170 4.280 ;
        RECT 813.010 4.000 814.010 4.280 ;
        RECT 814.850 4.000 815.850 4.280 ;
        RECT 816.690 4.000 817.690 4.280 ;
        RECT 818.530 4.000 819.530 4.280 ;
        RECT 820.370 4.000 821.370 4.280 ;
        RECT 822.210 4.000 823.210 4.280 ;
        RECT 824.050 4.000 825.050 4.280 ;
        RECT 825.890 4.000 826.890 4.280 ;
        RECT 827.730 4.000 828.730 4.280 ;
        RECT 829.570 4.000 830.570 4.280 ;
        RECT 831.410 4.000 832.410 4.280 ;
        RECT 833.250 4.000 834.250 4.280 ;
        RECT 835.090 4.000 836.090 4.280 ;
        RECT 836.930 4.000 837.930 4.280 ;
        RECT 838.770 4.000 839.770 4.280 ;
        RECT 840.610 4.000 841.610 4.280 ;
        RECT 842.450 4.000 843.450 4.280 ;
        RECT 844.290 4.000 845.290 4.280 ;
        RECT 846.130 4.000 847.130 4.280 ;
        RECT 847.970 4.000 848.970 4.280 ;
        RECT 849.810 4.000 850.810 4.280 ;
        RECT 851.650 4.000 852.650 4.280 ;
        RECT 853.490 4.000 854.490 4.280 ;
        RECT 855.330 4.000 856.330 4.280 ;
        RECT 857.170 4.000 858.170 4.280 ;
        RECT 859.010 4.000 860.010 4.280 ;
        RECT 860.850 4.000 861.850 4.280 ;
        RECT 862.690 4.000 863.690 4.280 ;
        RECT 864.530 4.000 865.530 4.280 ;
        RECT 866.370 4.000 867.370 4.280 ;
        RECT 868.210 4.000 869.210 4.280 ;
        RECT 870.050 4.000 871.050 4.280 ;
        RECT 871.890 4.000 872.890 4.280 ;
        RECT 873.730 4.000 874.730 4.280 ;
        RECT 875.570 4.000 876.570 4.280 ;
        RECT 877.410 4.000 878.410 4.280 ;
        RECT 879.250 4.000 880.250 4.280 ;
        RECT 881.090 4.000 882.090 4.280 ;
        RECT 882.930 4.000 883.930 4.280 ;
        RECT 884.770 4.000 885.770 4.280 ;
        RECT 886.610 4.000 887.610 4.280 ;
        RECT 888.450 4.000 889.450 4.280 ;
        RECT 890.290 4.000 891.290 4.280 ;
        RECT 892.130 4.000 893.130 4.280 ;
        RECT 893.970 4.000 894.970 4.280 ;
        RECT 895.810 4.000 896.810 4.280 ;
        RECT 897.650 4.000 898.650 4.280 ;
      LAYER met3 ;
        RECT 4.000 300.920 896.000 587.685 ;
        RECT 4.400 299.520 895.600 300.920 ;
        RECT 4.000 10.715 896.000 299.520 ;
      LAYER met4 ;
        RECT 8.150 18.110 20.640 430.945 ;
        RECT 23.040 18.110 23.940 430.945 ;
        RECT 26.340 18.110 27.240 430.945 ;
        RECT 29.640 18.110 30.540 430.945 ;
        RECT 32.940 18.110 97.440 430.945 ;
        RECT 99.840 18.110 100.740 430.945 ;
        RECT 103.140 18.110 104.040 430.945 ;
        RECT 106.440 18.110 107.340 430.945 ;
        RECT 109.740 18.110 174.240 430.945 ;
        RECT 176.640 18.110 177.540 430.945 ;
        RECT 179.940 18.110 180.840 430.945 ;
        RECT 183.240 18.110 184.140 430.945 ;
        RECT 186.540 18.110 251.040 430.945 ;
        RECT 253.440 18.110 254.340 430.945 ;
        RECT 256.740 18.110 257.640 430.945 ;
        RECT 260.040 18.110 260.940 430.945 ;
        RECT 263.340 18.110 327.840 430.945 ;
        RECT 330.240 18.110 331.140 430.945 ;
        RECT 333.540 18.110 334.440 430.945 ;
        RECT 336.840 18.110 337.740 430.945 ;
        RECT 340.140 18.110 404.640 430.945 ;
        RECT 407.040 18.110 407.940 430.945 ;
        RECT 410.340 18.110 411.240 430.945 ;
        RECT 413.640 18.110 414.540 430.945 ;
        RECT 416.940 18.110 481.440 430.945 ;
        RECT 483.840 18.110 484.740 430.945 ;
        RECT 487.140 18.110 488.040 430.945 ;
        RECT 490.440 18.110 491.340 430.945 ;
        RECT 493.740 18.110 558.240 430.945 ;
        RECT 560.640 18.110 561.540 430.945 ;
        RECT 563.940 18.110 564.840 430.945 ;
        RECT 567.240 18.110 568.140 430.945 ;
        RECT 570.540 18.110 635.040 430.945 ;
        RECT 637.440 18.110 638.185 430.945 ;
      LAYER met5 ;
        RECT 7.940 17.900 553.260 19.500 ;
  END
END user_proj
END LIBRARY

