magic
tech sky130A
magscale 1 2
timestamp 1624875440
<< obsli1 >>
rect 1104 1105 296884 295409
<< obsm1 >>
rect 290 960 297698 295440
<< metal2 >>
rect 1214 297200 1270 298000
rect 3698 297200 3754 298000
rect 6274 297200 6330 298000
rect 8850 297200 8906 298000
rect 11426 297200 11482 298000
rect 14002 297200 14058 298000
rect 16578 297200 16634 298000
rect 19154 297200 19210 298000
rect 21730 297200 21786 298000
rect 24306 297200 24362 298000
rect 26882 297200 26938 298000
rect 29458 297200 29514 298000
rect 32034 297200 32090 298000
rect 34518 297200 34574 298000
rect 37094 297200 37150 298000
rect 39670 297200 39726 298000
rect 42246 297200 42302 298000
rect 44822 297200 44878 298000
rect 47398 297200 47454 298000
rect 49974 297200 50030 298000
rect 52550 297200 52606 298000
rect 55126 297200 55182 298000
rect 57702 297200 57758 298000
rect 60278 297200 60334 298000
rect 62854 297200 62910 298000
rect 65430 297200 65486 298000
rect 67914 297200 67970 298000
rect 70490 297200 70546 298000
rect 73066 297200 73122 298000
rect 75642 297200 75698 298000
rect 78218 297200 78274 298000
rect 80794 297200 80850 298000
rect 83370 297200 83426 298000
rect 85946 297200 86002 298000
rect 88522 297200 88578 298000
rect 91098 297200 91154 298000
rect 93674 297200 93730 298000
rect 96250 297200 96306 298000
rect 98826 297200 98882 298000
rect 101310 297200 101366 298000
rect 103886 297200 103942 298000
rect 106462 297200 106518 298000
rect 109038 297200 109094 298000
rect 111614 297200 111670 298000
rect 114190 297200 114246 298000
rect 116766 297200 116822 298000
rect 119342 297200 119398 298000
rect 121918 297200 121974 298000
rect 124494 297200 124550 298000
rect 127070 297200 127126 298000
rect 129646 297200 129702 298000
rect 132222 297200 132278 298000
rect 134706 297200 134762 298000
rect 137282 297200 137338 298000
rect 139858 297200 139914 298000
rect 142434 297200 142490 298000
rect 145010 297200 145066 298000
rect 147586 297200 147642 298000
rect 150162 297200 150218 298000
rect 152738 297200 152794 298000
rect 155314 297200 155370 298000
rect 157890 297200 157946 298000
rect 160466 297200 160522 298000
rect 163042 297200 163098 298000
rect 165618 297200 165674 298000
rect 168102 297200 168158 298000
rect 170678 297200 170734 298000
rect 173254 297200 173310 298000
rect 175830 297200 175886 298000
rect 178406 297200 178462 298000
rect 180982 297200 181038 298000
rect 183558 297200 183614 298000
rect 186134 297200 186190 298000
rect 188710 297200 188766 298000
rect 191286 297200 191342 298000
rect 193862 297200 193918 298000
rect 196438 297200 196494 298000
rect 199014 297200 199070 298000
rect 201498 297200 201554 298000
rect 204074 297200 204130 298000
rect 206650 297200 206706 298000
rect 209226 297200 209282 298000
rect 211802 297200 211858 298000
rect 214378 297200 214434 298000
rect 216954 297200 217010 298000
rect 219530 297200 219586 298000
rect 222106 297200 222162 298000
rect 224682 297200 224738 298000
rect 227258 297200 227314 298000
rect 229834 297200 229890 298000
rect 232410 297200 232466 298000
rect 234894 297200 234950 298000
rect 237470 297200 237526 298000
rect 240046 297200 240102 298000
rect 242622 297200 242678 298000
rect 245198 297200 245254 298000
rect 247774 297200 247830 298000
rect 250350 297200 250406 298000
rect 252926 297200 252982 298000
rect 255502 297200 255558 298000
rect 258078 297200 258134 298000
rect 260654 297200 260710 298000
rect 263230 297200 263286 298000
rect 265806 297200 265862 298000
rect 268290 297200 268346 298000
rect 270866 297200 270922 298000
rect 273442 297200 273498 298000
rect 276018 297200 276074 298000
rect 278594 297200 278650 298000
rect 281170 297200 281226 298000
rect 283746 297200 283802 298000
rect 286322 297200 286378 298000
rect 288898 297200 288954 298000
rect 291474 297200 291530 298000
rect 294050 297200 294106 298000
rect 296626 297200 296682 298000
rect 294 0 350 800
rect 846 0 902 800
rect 1490 0 1546 800
rect 2042 0 2098 800
rect 2686 0 2742 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5722 0 5778 800
rect 6274 0 6330 800
rect 6918 0 6974 800
rect 7562 0 7618 800
rect 8114 0 8170 800
rect 8758 0 8814 800
rect 9310 0 9366 800
rect 9954 0 10010 800
rect 10598 0 10654 800
rect 11150 0 11206 800
rect 11794 0 11850 800
rect 12346 0 12402 800
rect 12990 0 13046 800
rect 13634 0 13690 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15382 0 15438 800
rect 16026 0 16082 800
rect 16670 0 16726 800
rect 17222 0 17278 800
rect 17866 0 17922 800
rect 18418 0 18474 800
rect 19062 0 19118 800
rect 19706 0 19762 800
rect 20258 0 20314 800
rect 20902 0 20958 800
rect 21454 0 21510 800
rect 22098 0 22154 800
rect 22742 0 22798 800
rect 23294 0 23350 800
rect 23938 0 23994 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26330 0 26386 800
rect 26974 0 27030 800
rect 27526 0 27582 800
rect 28170 0 28226 800
rect 28814 0 28870 800
rect 29366 0 29422 800
rect 30010 0 30066 800
rect 30562 0 30618 800
rect 31206 0 31262 800
rect 31850 0 31906 800
rect 32402 0 32458 800
rect 33046 0 33102 800
rect 33598 0 33654 800
rect 34242 0 34298 800
rect 34886 0 34942 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36634 0 36690 800
rect 37278 0 37334 800
rect 37830 0 37886 800
rect 38474 0 38530 800
rect 39118 0 39174 800
rect 39670 0 39726 800
rect 40314 0 40370 800
rect 40866 0 40922 800
rect 41510 0 41566 800
rect 42154 0 42210 800
rect 42706 0 42762 800
rect 43350 0 43406 800
rect 43902 0 43958 800
rect 44546 0 44602 800
rect 45190 0 45246 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 46938 0 46994 800
rect 47582 0 47638 800
rect 48226 0 48282 800
rect 48778 0 48834 800
rect 49422 0 49478 800
rect 49974 0 50030 800
rect 50618 0 50674 800
rect 51262 0 51318 800
rect 51814 0 51870 800
rect 52458 0 52514 800
rect 53010 0 53066 800
rect 53654 0 53710 800
rect 54298 0 54354 800
rect 54850 0 54906 800
rect 55494 0 55550 800
rect 56046 0 56102 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57886 0 57942 800
rect 58530 0 58586 800
rect 59082 0 59138 800
rect 59726 0 59782 800
rect 60370 0 60426 800
rect 60922 0 60978 800
rect 61566 0 61622 800
rect 62118 0 62174 800
rect 62762 0 62818 800
rect 63406 0 63462 800
rect 63958 0 64014 800
rect 64602 0 64658 800
rect 65154 0 65210 800
rect 65798 0 65854 800
rect 66442 0 66498 800
rect 66994 0 67050 800
rect 67638 0 67694 800
rect 68190 0 68246 800
rect 68834 0 68890 800
rect 69478 0 69534 800
rect 70030 0 70086 800
rect 70674 0 70730 800
rect 71226 0 71282 800
rect 71870 0 71926 800
rect 72514 0 72570 800
rect 73066 0 73122 800
rect 73710 0 73766 800
rect 74262 0 74318 800
rect 74906 0 74962 800
rect 75458 0 75514 800
rect 76102 0 76158 800
rect 76746 0 76802 800
rect 77298 0 77354 800
rect 77942 0 77998 800
rect 78494 0 78550 800
rect 79138 0 79194 800
rect 79782 0 79838 800
rect 80334 0 80390 800
rect 80978 0 81034 800
rect 81530 0 81586 800
rect 82174 0 82230 800
rect 82818 0 82874 800
rect 83370 0 83426 800
rect 84014 0 84070 800
rect 84566 0 84622 800
rect 85210 0 85266 800
rect 85854 0 85910 800
rect 86406 0 86462 800
rect 87050 0 87106 800
rect 87602 0 87658 800
rect 88246 0 88302 800
rect 88890 0 88946 800
rect 89442 0 89498 800
rect 90086 0 90142 800
rect 90638 0 90694 800
rect 91282 0 91338 800
rect 91926 0 91982 800
rect 92478 0 92534 800
rect 93122 0 93178 800
rect 93674 0 93730 800
rect 94318 0 94374 800
rect 94962 0 95018 800
rect 95514 0 95570 800
rect 96158 0 96214 800
rect 96710 0 96766 800
rect 97354 0 97410 800
rect 97998 0 98054 800
rect 98550 0 98606 800
rect 99194 0 99250 800
rect 99746 0 99802 800
rect 100390 0 100446 800
rect 101034 0 101090 800
rect 101586 0 101642 800
rect 102230 0 102286 800
rect 102782 0 102838 800
rect 103426 0 103482 800
rect 104070 0 104126 800
rect 104622 0 104678 800
rect 105266 0 105322 800
rect 105818 0 105874 800
rect 106462 0 106518 800
rect 107106 0 107162 800
rect 107658 0 107714 800
rect 108302 0 108358 800
rect 108854 0 108910 800
rect 109498 0 109554 800
rect 110142 0 110198 800
rect 110694 0 110750 800
rect 111338 0 111394 800
rect 111890 0 111946 800
rect 112534 0 112590 800
rect 113086 0 113142 800
rect 113730 0 113786 800
rect 114374 0 114430 800
rect 114926 0 114982 800
rect 115570 0 115626 800
rect 116122 0 116178 800
rect 116766 0 116822 800
rect 117410 0 117466 800
rect 117962 0 118018 800
rect 118606 0 118662 800
rect 119158 0 119214 800
rect 119802 0 119858 800
rect 120446 0 120502 800
rect 120998 0 121054 800
rect 121642 0 121698 800
rect 122194 0 122250 800
rect 122838 0 122894 800
rect 123482 0 123538 800
rect 124034 0 124090 800
rect 124678 0 124734 800
rect 125230 0 125286 800
rect 125874 0 125930 800
rect 126518 0 126574 800
rect 127070 0 127126 800
rect 127714 0 127770 800
rect 128266 0 128322 800
rect 128910 0 128966 800
rect 129554 0 129610 800
rect 130106 0 130162 800
rect 130750 0 130806 800
rect 131302 0 131358 800
rect 131946 0 132002 800
rect 132590 0 132646 800
rect 133142 0 133198 800
rect 133786 0 133842 800
rect 134338 0 134394 800
rect 134982 0 135038 800
rect 135626 0 135682 800
rect 136178 0 136234 800
rect 136822 0 136878 800
rect 137374 0 137430 800
rect 138018 0 138074 800
rect 138662 0 138718 800
rect 139214 0 139270 800
rect 139858 0 139914 800
rect 140410 0 140466 800
rect 141054 0 141110 800
rect 141698 0 141754 800
rect 142250 0 142306 800
rect 142894 0 142950 800
rect 143446 0 143502 800
rect 144090 0 144146 800
rect 144734 0 144790 800
rect 145286 0 145342 800
rect 145930 0 145986 800
rect 146482 0 146538 800
rect 147126 0 147182 800
rect 147770 0 147826 800
rect 148322 0 148378 800
rect 148966 0 149022 800
rect 149518 0 149574 800
rect 150162 0 150218 800
rect 150714 0 150770 800
rect 151358 0 151414 800
rect 152002 0 152058 800
rect 152554 0 152610 800
rect 153198 0 153254 800
rect 153750 0 153806 800
rect 154394 0 154450 800
rect 155038 0 155094 800
rect 155590 0 155646 800
rect 156234 0 156290 800
rect 156786 0 156842 800
rect 157430 0 157486 800
rect 158074 0 158130 800
rect 158626 0 158682 800
rect 159270 0 159326 800
rect 159822 0 159878 800
rect 160466 0 160522 800
rect 161110 0 161166 800
rect 161662 0 161718 800
rect 162306 0 162362 800
rect 162858 0 162914 800
rect 163502 0 163558 800
rect 164146 0 164202 800
rect 164698 0 164754 800
rect 165342 0 165398 800
rect 165894 0 165950 800
rect 166538 0 166594 800
rect 167182 0 167238 800
rect 167734 0 167790 800
rect 168378 0 168434 800
rect 168930 0 168986 800
rect 169574 0 169630 800
rect 170218 0 170274 800
rect 170770 0 170826 800
rect 171414 0 171470 800
rect 171966 0 172022 800
rect 172610 0 172666 800
rect 173254 0 173310 800
rect 173806 0 173862 800
rect 174450 0 174506 800
rect 175002 0 175058 800
rect 175646 0 175702 800
rect 176290 0 176346 800
rect 176842 0 176898 800
rect 177486 0 177542 800
rect 178038 0 178094 800
rect 178682 0 178738 800
rect 179326 0 179382 800
rect 179878 0 179934 800
rect 180522 0 180578 800
rect 181074 0 181130 800
rect 181718 0 181774 800
rect 182362 0 182418 800
rect 182914 0 182970 800
rect 183558 0 183614 800
rect 184110 0 184166 800
rect 184754 0 184810 800
rect 185398 0 185454 800
rect 185950 0 186006 800
rect 186594 0 186650 800
rect 187146 0 187202 800
rect 187790 0 187846 800
rect 188342 0 188398 800
rect 188986 0 189042 800
rect 189630 0 189686 800
rect 190182 0 190238 800
rect 190826 0 190882 800
rect 191378 0 191434 800
rect 192022 0 192078 800
rect 192666 0 192722 800
rect 193218 0 193274 800
rect 193862 0 193918 800
rect 194414 0 194470 800
rect 195058 0 195114 800
rect 195702 0 195758 800
rect 196254 0 196310 800
rect 196898 0 196954 800
rect 197450 0 197506 800
rect 198094 0 198150 800
rect 198738 0 198794 800
rect 199290 0 199346 800
rect 199934 0 199990 800
rect 200486 0 200542 800
rect 201130 0 201186 800
rect 201774 0 201830 800
rect 202326 0 202382 800
rect 202970 0 203026 800
rect 203522 0 203578 800
rect 204166 0 204222 800
rect 204810 0 204866 800
rect 205362 0 205418 800
rect 206006 0 206062 800
rect 206558 0 206614 800
rect 207202 0 207258 800
rect 207846 0 207902 800
rect 208398 0 208454 800
rect 209042 0 209098 800
rect 209594 0 209650 800
rect 210238 0 210294 800
rect 210882 0 210938 800
rect 211434 0 211490 800
rect 212078 0 212134 800
rect 212630 0 212686 800
rect 213274 0 213330 800
rect 213918 0 213974 800
rect 214470 0 214526 800
rect 215114 0 215170 800
rect 215666 0 215722 800
rect 216310 0 216366 800
rect 216954 0 217010 800
rect 217506 0 217562 800
rect 218150 0 218206 800
rect 218702 0 218758 800
rect 219346 0 219402 800
rect 219990 0 220046 800
rect 220542 0 220598 800
rect 221186 0 221242 800
rect 221738 0 221794 800
rect 222382 0 222438 800
rect 223026 0 223082 800
rect 223578 0 223634 800
rect 224222 0 224278 800
rect 224774 0 224830 800
rect 225418 0 225474 800
rect 225970 0 226026 800
rect 226614 0 226670 800
rect 227258 0 227314 800
rect 227810 0 227866 800
rect 228454 0 228510 800
rect 229006 0 229062 800
rect 229650 0 229706 800
rect 230294 0 230350 800
rect 230846 0 230902 800
rect 231490 0 231546 800
rect 232042 0 232098 800
rect 232686 0 232742 800
rect 233330 0 233386 800
rect 233882 0 233938 800
rect 234526 0 234582 800
rect 235078 0 235134 800
rect 235722 0 235778 800
rect 236366 0 236422 800
rect 236918 0 236974 800
rect 237562 0 237618 800
rect 238114 0 238170 800
rect 238758 0 238814 800
rect 239402 0 239458 800
rect 239954 0 240010 800
rect 240598 0 240654 800
rect 241150 0 241206 800
rect 241794 0 241850 800
rect 242438 0 242494 800
rect 242990 0 243046 800
rect 243634 0 243690 800
rect 244186 0 244242 800
rect 244830 0 244886 800
rect 245474 0 245530 800
rect 246026 0 246082 800
rect 246670 0 246726 800
rect 247222 0 247278 800
rect 247866 0 247922 800
rect 248510 0 248566 800
rect 249062 0 249118 800
rect 249706 0 249762 800
rect 250258 0 250314 800
rect 250902 0 250958 800
rect 251546 0 251602 800
rect 252098 0 252154 800
rect 252742 0 252798 800
rect 253294 0 253350 800
rect 253938 0 253994 800
rect 254582 0 254638 800
rect 255134 0 255190 800
rect 255778 0 255834 800
rect 256330 0 256386 800
rect 256974 0 257030 800
rect 257618 0 257674 800
rect 258170 0 258226 800
rect 258814 0 258870 800
rect 259366 0 259422 800
rect 260010 0 260066 800
rect 260654 0 260710 800
rect 261206 0 261262 800
rect 261850 0 261906 800
rect 262402 0 262458 800
rect 263046 0 263102 800
rect 263598 0 263654 800
rect 264242 0 264298 800
rect 264886 0 264942 800
rect 265438 0 265494 800
rect 266082 0 266138 800
rect 266634 0 266690 800
rect 267278 0 267334 800
rect 267922 0 267978 800
rect 268474 0 268530 800
rect 269118 0 269174 800
rect 269670 0 269726 800
rect 270314 0 270370 800
rect 270958 0 271014 800
rect 271510 0 271566 800
rect 272154 0 272210 800
rect 272706 0 272762 800
rect 273350 0 273406 800
rect 273994 0 274050 800
rect 274546 0 274602 800
rect 275190 0 275246 800
rect 275742 0 275798 800
rect 276386 0 276442 800
rect 277030 0 277086 800
rect 277582 0 277638 800
rect 278226 0 278282 800
rect 278778 0 278834 800
rect 279422 0 279478 800
rect 280066 0 280122 800
rect 280618 0 280674 800
rect 281262 0 281318 800
rect 281814 0 281870 800
rect 282458 0 282514 800
rect 283102 0 283158 800
rect 283654 0 283710 800
rect 284298 0 284354 800
rect 284850 0 284906 800
rect 285494 0 285550 800
rect 286138 0 286194 800
rect 286690 0 286746 800
rect 287334 0 287390 800
rect 287886 0 287942 800
rect 288530 0 288586 800
rect 289174 0 289230 800
rect 289726 0 289782 800
rect 290370 0 290426 800
rect 290922 0 290978 800
rect 291566 0 291622 800
rect 292210 0 292266 800
rect 292762 0 292818 800
rect 293406 0 293462 800
rect 293958 0 294014 800
rect 294602 0 294658 800
rect 295246 0 295302 800
rect 295798 0 295854 800
rect 296442 0 296498 800
rect 296994 0 297050 800
rect 297638 0 297694 800
<< obsm2 >>
rect 296 297144 1158 297200
rect 1326 297144 3642 297200
rect 3810 297144 6218 297200
rect 6386 297144 8794 297200
rect 8962 297144 11370 297200
rect 11538 297144 13946 297200
rect 14114 297144 16522 297200
rect 16690 297144 19098 297200
rect 19266 297144 21674 297200
rect 21842 297144 24250 297200
rect 24418 297144 26826 297200
rect 26994 297144 29402 297200
rect 29570 297144 31978 297200
rect 32146 297144 34462 297200
rect 34630 297144 37038 297200
rect 37206 297144 39614 297200
rect 39782 297144 42190 297200
rect 42358 297144 44766 297200
rect 44934 297144 47342 297200
rect 47510 297144 49918 297200
rect 50086 297144 52494 297200
rect 52662 297144 55070 297200
rect 55238 297144 57646 297200
rect 57814 297144 60222 297200
rect 60390 297144 62798 297200
rect 62966 297144 65374 297200
rect 65542 297144 67858 297200
rect 68026 297144 70434 297200
rect 70602 297144 73010 297200
rect 73178 297144 75586 297200
rect 75754 297144 78162 297200
rect 78330 297144 80738 297200
rect 80906 297144 83314 297200
rect 83482 297144 85890 297200
rect 86058 297144 88466 297200
rect 88634 297144 91042 297200
rect 91210 297144 93618 297200
rect 93786 297144 96194 297200
rect 96362 297144 98770 297200
rect 98938 297144 101254 297200
rect 101422 297144 103830 297200
rect 103998 297144 106406 297200
rect 106574 297144 108982 297200
rect 109150 297144 111558 297200
rect 111726 297144 114134 297200
rect 114302 297144 116710 297200
rect 116878 297144 119286 297200
rect 119454 297144 121862 297200
rect 122030 297144 124438 297200
rect 124606 297144 127014 297200
rect 127182 297144 129590 297200
rect 129758 297144 132166 297200
rect 132334 297144 134650 297200
rect 134818 297144 137226 297200
rect 137394 297144 139802 297200
rect 139970 297144 142378 297200
rect 142546 297144 144954 297200
rect 145122 297144 147530 297200
rect 147698 297144 150106 297200
rect 150274 297144 152682 297200
rect 152850 297144 155258 297200
rect 155426 297144 157834 297200
rect 158002 297144 160410 297200
rect 160578 297144 162986 297200
rect 163154 297144 165562 297200
rect 165730 297144 168046 297200
rect 168214 297144 170622 297200
rect 170790 297144 173198 297200
rect 173366 297144 175774 297200
rect 175942 297144 178350 297200
rect 178518 297144 180926 297200
rect 181094 297144 183502 297200
rect 183670 297144 186078 297200
rect 186246 297144 188654 297200
rect 188822 297144 191230 297200
rect 191398 297144 193806 297200
rect 193974 297144 196382 297200
rect 196550 297144 198958 297200
rect 199126 297144 201442 297200
rect 201610 297144 204018 297200
rect 204186 297144 206594 297200
rect 206762 297144 209170 297200
rect 209338 297144 211746 297200
rect 211914 297144 214322 297200
rect 214490 297144 216898 297200
rect 217066 297144 219474 297200
rect 219642 297144 222050 297200
rect 222218 297144 224626 297200
rect 224794 297144 227202 297200
rect 227370 297144 229778 297200
rect 229946 297144 232354 297200
rect 232522 297144 234838 297200
rect 235006 297144 237414 297200
rect 237582 297144 239990 297200
rect 240158 297144 242566 297200
rect 242734 297144 245142 297200
rect 245310 297144 247718 297200
rect 247886 297144 250294 297200
rect 250462 297144 252870 297200
rect 253038 297144 255446 297200
rect 255614 297144 258022 297200
rect 258190 297144 260598 297200
rect 260766 297144 263174 297200
rect 263342 297144 265750 297200
rect 265918 297144 268234 297200
rect 268402 297144 270810 297200
rect 270978 297144 273386 297200
rect 273554 297144 275962 297200
rect 276130 297144 278538 297200
rect 278706 297144 281114 297200
rect 281282 297144 283690 297200
rect 283858 297144 286266 297200
rect 286434 297144 288842 297200
rect 289010 297144 291418 297200
rect 291586 297144 293994 297200
rect 294162 297144 296570 297200
rect 296738 297144 297692 297200
rect 296 856 297692 297144
rect 406 800 790 856
rect 958 800 1434 856
rect 1602 800 1986 856
rect 2154 800 2630 856
rect 2798 800 3182 856
rect 3350 800 3826 856
rect 3994 800 4470 856
rect 4638 800 5022 856
rect 5190 800 5666 856
rect 5834 800 6218 856
rect 6386 800 6862 856
rect 7030 800 7506 856
rect 7674 800 8058 856
rect 8226 800 8702 856
rect 8870 800 9254 856
rect 9422 800 9898 856
rect 10066 800 10542 856
rect 10710 800 11094 856
rect 11262 800 11738 856
rect 11906 800 12290 856
rect 12458 800 12934 856
rect 13102 800 13578 856
rect 13746 800 14130 856
rect 14298 800 14774 856
rect 14942 800 15326 856
rect 15494 800 15970 856
rect 16138 800 16614 856
rect 16782 800 17166 856
rect 17334 800 17810 856
rect 17978 800 18362 856
rect 18530 800 19006 856
rect 19174 800 19650 856
rect 19818 800 20202 856
rect 20370 800 20846 856
rect 21014 800 21398 856
rect 21566 800 22042 856
rect 22210 800 22686 856
rect 22854 800 23238 856
rect 23406 800 23882 856
rect 24050 800 24434 856
rect 24602 800 25078 856
rect 25246 800 25722 856
rect 25890 800 26274 856
rect 26442 800 26918 856
rect 27086 800 27470 856
rect 27638 800 28114 856
rect 28282 800 28758 856
rect 28926 800 29310 856
rect 29478 800 29954 856
rect 30122 800 30506 856
rect 30674 800 31150 856
rect 31318 800 31794 856
rect 31962 800 32346 856
rect 32514 800 32990 856
rect 33158 800 33542 856
rect 33710 800 34186 856
rect 34354 800 34830 856
rect 34998 800 35382 856
rect 35550 800 36026 856
rect 36194 800 36578 856
rect 36746 800 37222 856
rect 37390 800 37774 856
rect 37942 800 38418 856
rect 38586 800 39062 856
rect 39230 800 39614 856
rect 39782 800 40258 856
rect 40426 800 40810 856
rect 40978 800 41454 856
rect 41622 800 42098 856
rect 42266 800 42650 856
rect 42818 800 43294 856
rect 43462 800 43846 856
rect 44014 800 44490 856
rect 44658 800 45134 856
rect 45302 800 45686 856
rect 45854 800 46330 856
rect 46498 800 46882 856
rect 47050 800 47526 856
rect 47694 800 48170 856
rect 48338 800 48722 856
rect 48890 800 49366 856
rect 49534 800 49918 856
rect 50086 800 50562 856
rect 50730 800 51206 856
rect 51374 800 51758 856
rect 51926 800 52402 856
rect 52570 800 52954 856
rect 53122 800 53598 856
rect 53766 800 54242 856
rect 54410 800 54794 856
rect 54962 800 55438 856
rect 55606 800 55990 856
rect 56158 800 56634 856
rect 56802 800 57278 856
rect 57446 800 57830 856
rect 57998 800 58474 856
rect 58642 800 59026 856
rect 59194 800 59670 856
rect 59838 800 60314 856
rect 60482 800 60866 856
rect 61034 800 61510 856
rect 61678 800 62062 856
rect 62230 800 62706 856
rect 62874 800 63350 856
rect 63518 800 63902 856
rect 64070 800 64546 856
rect 64714 800 65098 856
rect 65266 800 65742 856
rect 65910 800 66386 856
rect 66554 800 66938 856
rect 67106 800 67582 856
rect 67750 800 68134 856
rect 68302 800 68778 856
rect 68946 800 69422 856
rect 69590 800 69974 856
rect 70142 800 70618 856
rect 70786 800 71170 856
rect 71338 800 71814 856
rect 71982 800 72458 856
rect 72626 800 73010 856
rect 73178 800 73654 856
rect 73822 800 74206 856
rect 74374 800 74850 856
rect 75018 800 75402 856
rect 75570 800 76046 856
rect 76214 800 76690 856
rect 76858 800 77242 856
rect 77410 800 77886 856
rect 78054 800 78438 856
rect 78606 800 79082 856
rect 79250 800 79726 856
rect 79894 800 80278 856
rect 80446 800 80922 856
rect 81090 800 81474 856
rect 81642 800 82118 856
rect 82286 800 82762 856
rect 82930 800 83314 856
rect 83482 800 83958 856
rect 84126 800 84510 856
rect 84678 800 85154 856
rect 85322 800 85798 856
rect 85966 800 86350 856
rect 86518 800 86994 856
rect 87162 800 87546 856
rect 87714 800 88190 856
rect 88358 800 88834 856
rect 89002 800 89386 856
rect 89554 800 90030 856
rect 90198 800 90582 856
rect 90750 800 91226 856
rect 91394 800 91870 856
rect 92038 800 92422 856
rect 92590 800 93066 856
rect 93234 800 93618 856
rect 93786 800 94262 856
rect 94430 800 94906 856
rect 95074 800 95458 856
rect 95626 800 96102 856
rect 96270 800 96654 856
rect 96822 800 97298 856
rect 97466 800 97942 856
rect 98110 800 98494 856
rect 98662 800 99138 856
rect 99306 800 99690 856
rect 99858 800 100334 856
rect 100502 800 100978 856
rect 101146 800 101530 856
rect 101698 800 102174 856
rect 102342 800 102726 856
rect 102894 800 103370 856
rect 103538 800 104014 856
rect 104182 800 104566 856
rect 104734 800 105210 856
rect 105378 800 105762 856
rect 105930 800 106406 856
rect 106574 800 107050 856
rect 107218 800 107602 856
rect 107770 800 108246 856
rect 108414 800 108798 856
rect 108966 800 109442 856
rect 109610 800 110086 856
rect 110254 800 110638 856
rect 110806 800 111282 856
rect 111450 800 111834 856
rect 112002 800 112478 856
rect 112646 800 113030 856
rect 113198 800 113674 856
rect 113842 800 114318 856
rect 114486 800 114870 856
rect 115038 800 115514 856
rect 115682 800 116066 856
rect 116234 800 116710 856
rect 116878 800 117354 856
rect 117522 800 117906 856
rect 118074 800 118550 856
rect 118718 800 119102 856
rect 119270 800 119746 856
rect 119914 800 120390 856
rect 120558 800 120942 856
rect 121110 800 121586 856
rect 121754 800 122138 856
rect 122306 800 122782 856
rect 122950 800 123426 856
rect 123594 800 123978 856
rect 124146 800 124622 856
rect 124790 800 125174 856
rect 125342 800 125818 856
rect 125986 800 126462 856
rect 126630 800 127014 856
rect 127182 800 127658 856
rect 127826 800 128210 856
rect 128378 800 128854 856
rect 129022 800 129498 856
rect 129666 800 130050 856
rect 130218 800 130694 856
rect 130862 800 131246 856
rect 131414 800 131890 856
rect 132058 800 132534 856
rect 132702 800 133086 856
rect 133254 800 133730 856
rect 133898 800 134282 856
rect 134450 800 134926 856
rect 135094 800 135570 856
rect 135738 800 136122 856
rect 136290 800 136766 856
rect 136934 800 137318 856
rect 137486 800 137962 856
rect 138130 800 138606 856
rect 138774 800 139158 856
rect 139326 800 139802 856
rect 139970 800 140354 856
rect 140522 800 140998 856
rect 141166 800 141642 856
rect 141810 800 142194 856
rect 142362 800 142838 856
rect 143006 800 143390 856
rect 143558 800 144034 856
rect 144202 800 144678 856
rect 144846 800 145230 856
rect 145398 800 145874 856
rect 146042 800 146426 856
rect 146594 800 147070 856
rect 147238 800 147714 856
rect 147882 800 148266 856
rect 148434 800 148910 856
rect 149078 800 149462 856
rect 149630 800 150106 856
rect 150274 800 150658 856
rect 150826 800 151302 856
rect 151470 800 151946 856
rect 152114 800 152498 856
rect 152666 800 153142 856
rect 153310 800 153694 856
rect 153862 800 154338 856
rect 154506 800 154982 856
rect 155150 800 155534 856
rect 155702 800 156178 856
rect 156346 800 156730 856
rect 156898 800 157374 856
rect 157542 800 158018 856
rect 158186 800 158570 856
rect 158738 800 159214 856
rect 159382 800 159766 856
rect 159934 800 160410 856
rect 160578 800 161054 856
rect 161222 800 161606 856
rect 161774 800 162250 856
rect 162418 800 162802 856
rect 162970 800 163446 856
rect 163614 800 164090 856
rect 164258 800 164642 856
rect 164810 800 165286 856
rect 165454 800 165838 856
rect 166006 800 166482 856
rect 166650 800 167126 856
rect 167294 800 167678 856
rect 167846 800 168322 856
rect 168490 800 168874 856
rect 169042 800 169518 856
rect 169686 800 170162 856
rect 170330 800 170714 856
rect 170882 800 171358 856
rect 171526 800 171910 856
rect 172078 800 172554 856
rect 172722 800 173198 856
rect 173366 800 173750 856
rect 173918 800 174394 856
rect 174562 800 174946 856
rect 175114 800 175590 856
rect 175758 800 176234 856
rect 176402 800 176786 856
rect 176954 800 177430 856
rect 177598 800 177982 856
rect 178150 800 178626 856
rect 178794 800 179270 856
rect 179438 800 179822 856
rect 179990 800 180466 856
rect 180634 800 181018 856
rect 181186 800 181662 856
rect 181830 800 182306 856
rect 182474 800 182858 856
rect 183026 800 183502 856
rect 183670 800 184054 856
rect 184222 800 184698 856
rect 184866 800 185342 856
rect 185510 800 185894 856
rect 186062 800 186538 856
rect 186706 800 187090 856
rect 187258 800 187734 856
rect 187902 800 188286 856
rect 188454 800 188930 856
rect 189098 800 189574 856
rect 189742 800 190126 856
rect 190294 800 190770 856
rect 190938 800 191322 856
rect 191490 800 191966 856
rect 192134 800 192610 856
rect 192778 800 193162 856
rect 193330 800 193806 856
rect 193974 800 194358 856
rect 194526 800 195002 856
rect 195170 800 195646 856
rect 195814 800 196198 856
rect 196366 800 196842 856
rect 197010 800 197394 856
rect 197562 800 198038 856
rect 198206 800 198682 856
rect 198850 800 199234 856
rect 199402 800 199878 856
rect 200046 800 200430 856
rect 200598 800 201074 856
rect 201242 800 201718 856
rect 201886 800 202270 856
rect 202438 800 202914 856
rect 203082 800 203466 856
rect 203634 800 204110 856
rect 204278 800 204754 856
rect 204922 800 205306 856
rect 205474 800 205950 856
rect 206118 800 206502 856
rect 206670 800 207146 856
rect 207314 800 207790 856
rect 207958 800 208342 856
rect 208510 800 208986 856
rect 209154 800 209538 856
rect 209706 800 210182 856
rect 210350 800 210826 856
rect 210994 800 211378 856
rect 211546 800 212022 856
rect 212190 800 212574 856
rect 212742 800 213218 856
rect 213386 800 213862 856
rect 214030 800 214414 856
rect 214582 800 215058 856
rect 215226 800 215610 856
rect 215778 800 216254 856
rect 216422 800 216898 856
rect 217066 800 217450 856
rect 217618 800 218094 856
rect 218262 800 218646 856
rect 218814 800 219290 856
rect 219458 800 219934 856
rect 220102 800 220486 856
rect 220654 800 221130 856
rect 221298 800 221682 856
rect 221850 800 222326 856
rect 222494 800 222970 856
rect 223138 800 223522 856
rect 223690 800 224166 856
rect 224334 800 224718 856
rect 224886 800 225362 856
rect 225530 800 225914 856
rect 226082 800 226558 856
rect 226726 800 227202 856
rect 227370 800 227754 856
rect 227922 800 228398 856
rect 228566 800 228950 856
rect 229118 800 229594 856
rect 229762 800 230238 856
rect 230406 800 230790 856
rect 230958 800 231434 856
rect 231602 800 231986 856
rect 232154 800 232630 856
rect 232798 800 233274 856
rect 233442 800 233826 856
rect 233994 800 234470 856
rect 234638 800 235022 856
rect 235190 800 235666 856
rect 235834 800 236310 856
rect 236478 800 236862 856
rect 237030 800 237506 856
rect 237674 800 238058 856
rect 238226 800 238702 856
rect 238870 800 239346 856
rect 239514 800 239898 856
rect 240066 800 240542 856
rect 240710 800 241094 856
rect 241262 800 241738 856
rect 241906 800 242382 856
rect 242550 800 242934 856
rect 243102 800 243578 856
rect 243746 800 244130 856
rect 244298 800 244774 856
rect 244942 800 245418 856
rect 245586 800 245970 856
rect 246138 800 246614 856
rect 246782 800 247166 856
rect 247334 800 247810 856
rect 247978 800 248454 856
rect 248622 800 249006 856
rect 249174 800 249650 856
rect 249818 800 250202 856
rect 250370 800 250846 856
rect 251014 800 251490 856
rect 251658 800 252042 856
rect 252210 800 252686 856
rect 252854 800 253238 856
rect 253406 800 253882 856
rect 254050 800 254526 856
rect 254694 800 255078 856
rect 255246 800 255722 856
rect 255890 800 256274 856
rect 256442 800 256918 856
rect 257086 800 257562 856
rect 257730 800 258114 856
rect 258282 800 258758 856
rect 258926 800 259310 856
rect 259478 800 259954 856
rect 260122 800 260598 856
rect 260766 800 261150 856
rect 261318 800 261794 856
rect 261962 800 262346 856
rect 262514 800 262990 856
rect 263158 800 263542 856
rect 263710 800 264186 856
rect 264354 800 264830 856
rect 264998 800 265382 856
rect 265550 800 266026 856
rect 266194 800 266578 856
rect 266746 800 267222 856
rect 267390 800 267866 856
rect 268034 800 268418 856
rect 268586 800 269062 856
rect 269230 800 269614 856
rect 269782 800 270258 856
rect 270426 800 270902 856
rect 271070 800 271454 856
rect 271622 800 272098 856
rect 272266 800 272650 856
rect 272818 800 273294 856
rect 273462 800 273938 856
rect 274106 800 274490 856
rect 274658 800 275134 856
rect 275302 800 275686 856
rect 275854 800 276330 856
rect 276498 800 276974 856
rect 277142 800 277526 856
rect 277694 800 278170 856
rect 278338 800 278722 856
rect 278890 800 279366 856
rect 279534 800 280010 856
rect 280178 800 280562 856
rect 280730 800 281206 856
rect 281374 800 281758 856
rect 281926 800 282402 856
rect 282570 800 283046 856
rect 283214 800 283598 856
rect 283766 800 284242 856
rect 284410 800 284794 856
rect 284962 800 285438 856
rect 285606 800 286082 856
rect 286250 800 286634 856
rect 286802 800 287278 856
rect 287446 800 287830 856
rect 287998 800 288474 856
rect 288642 800 289118 856
rect 289286 800 289670 856
rect 289838 800 290314 856
rect 290482 800 290866 856
rect 291034 800 291510 856
rect 291678 800 292154 856
rect 292322 800 292706 856
rect 292874 800 293350 856
rect 293518 800 293902 856
rect 294070 800 294546 856
rect 294714 800 295190 856
rect 295358 800 295742 856
rect 295910 800 296386 856
rect 296554 800 296938 856
rect 297106 800 297582 856
<< metal3 >>
rect 0 148928 800 149048
<< obsm3 >>
rect 800 149128 296687 295425
rect 880 148848 296687 149128
rect 800 1395 296687 148848
<< metal4 >>
rect 4208 2128 4528 295440
rect 4868 2176 5188 295392
rect 5528 2176 5848 295392
rect 6188 2176 6508 295392
rect 19568 2128 19888 295440
rect 20228 2176 20548 295392
rect 20888 2176 21208 295392
rect 21548 2176 21868 295392
rect 34928 2128 35248 295440
rect 35588 2176 35908 295392
rect 36248 2176 36568 295392
rect 36908 2176 37228 295392
rect 50288 2128 50608 295440
rect 50948 2176 51268 295392
rect 51608 2176 51928 295392
rect 52268 2176 52588 295392
rect 65648 2128 65968 295440
rect 66308 2176 66628 295392
rect 66968 2176 67288 295392
rect 67628 2176 67948 295392
rect 81008 2128 81328 295440
rect 81668 2176 81988 295392
rect 82328 2176 82648 295392
rect 82988 2176 83308 295392
rect 96368 2128 96688 295440
rect 97028 2176 97348 295392
rect 97688 2176 98008 295392
rect 98348 2176 98668 295392
rect 111728 2128 112048 295440
rect 112388 2176 112708 295392
rect 113048 2176 113368 295392
rect 113708 2176 114028 295392
rect 127088 2128 127408 295440
rect 127748 2176 128068 295392
rect 128408 2176 128728 295392
rect 129068 2176 129388 295392
rect 142448 2128 142768 295440
rect 143108 2176 143428 295392
rect 143768 2176 144088 295392
rect 144428 2176 144748 295392
rect 157808 2128 158128 295440
rect 158468 2176 158788 295392
rect 159128 2176 159448 295392
rect 159788 2176 160108 295392
rect 173168 2128 173488 295440
rect 173828 2176 174148 295392
rect 174488 2176 174808 295392
rect 175148 2176 175468 295392
rect 188528 2128 188848 295440
rect 189188 2176 189508 295392
rect 189848 2176 190168 295392
rect 190508 2176 190828 295392
rect 203888 2128 204208 295440
rect 204548 2176 204868 295392
rect 205208 2176 205528 295392
rect 205868 2176 206188 295392
rect 219248 2128 219568 295440
rect 219908 2176 220228 295392
rect 220568 2176 220888 295392
rect 221228 2176 221548 295392
rect 234608 2128 234928 295440
rect 235268 2176 235588 295392
rect 235928 2176 236248 295392
rect 236588 2176 236908 295392
rect 249968 2128 250288 295440
rect 250628 2176 250948 295392
rect 251288 2176 251608 295392
rect 251948 2176 252268 295392
rect 265328 2128 265648 295440
rect 265988 2176 266308 295392
rect 266648 2176 266968 295392
rect 267308 2176 267628 295392
rect 280688 2128 281008 295440
rect 281348 2176 281668 295392
rect 282008 2176 282328 295392
rect 282668 2176 282988 295392
rect 296048 2128 296368 295440
<< obsm4 >>
rect 4659 3163 4788 289645
rect 5268 3163 5448 289645
rect 5928 3163 6108 289645
rect 6588 3163 19488 289645
rect 19968 3163 20148 289645
rect 20628 3163 20808 289645
rect 21288 3163 21468 289645
rect 21948 3163 34848 289645
rect 35328 3163 35508 289645
rect 35988 3163 36168 289645
rect 36648 3163 36828 289645
rect 37308 3163 50208 289645
rect 50688 3163 50868 289645
rect 51348 3163 51528 289645
rect 52008 3163 52188 289645
rect 52668 3163 65568 289645
rect 66048 3163 66228 289645
rect 66708 3163 66888 289645
rect 67368 3163 67548 289645
rect 68028 3163 80928 289645
rect 81408 3163 81588 289645
rect 82068 3163 82248 289645
rect 82728 3163 82908 289645
rect 83388 3163 96288 289645
rect 96768 3163 96948 289645
rect 97428 3163 97608 289645
rect 98088 3163 98268 289645
rect 98748 3163 111648 289645
rect 112128 3163 112308 289645
rect 112788 3163 112968 289645
rect 113448 3163 113628 289645
rect 114108 3163 127008 289645
rect 127488 3163 127668 289645
rect 128148 3163 128328 289645
rect 128808 3163 128988 289645
rect 129468 3163 142368 289645
rect 142848 3163 143028 289645
rect 143508 3163 143688 289645
rect 144168 3163 144348 289645
rect 144828 3163 157728 289645
rect 158208 3163 158388 289645
rect 158868 3163 159048 289645
rect 159528 3163 159708 289645
rect 160188 3163 173088 289645
rect 173568 3163 173748 289645
rect 174228 3163 174408 289645
rect 174888 3163 175068 289645
rect 175548 3163 188448 289645
rect 188928 3163 189108 289645
rect 189588 3163 189768 289645
rect 190248 3163 190428 289645
rect 190908 3163 203808 289645
rect 204288 3163 204468 289645
rect 204948 3163 205128 289645
rect 205608 3163 205788 289645
rect 206268 3163 219168 289645
rect 219648 3163 219828 289645
rect 220308 3163 220488 289645
rect 220968 3163 221148 289645
rect 221628 3163 234528 289645
rect 235008 3163 235188 289645
rect 235668 3163 235848 289645
rect 236328 3163 236508 289645
rect 236988 3163 249888 289645
rect 250368 3163 250548 289645
rect 251028 3163 251208 289645
rect 251688 3163 251868 289645
rect 252348 3163 265248 289645
rect 265728 3163 265908 289645
rect 266388 3163 266568 289645
rect 267048 3163 267228 289645
rect 267708 3163 280608 289645
rect 281088 3163 281268 289645
rect 281748 3163 281928 289645
rect 282408 3163 282588 289645
rect 283068 3163 288269 289645
<< labels >>
rlabel metal2 s 1214 297200 1270 298000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 78218 297200 78274 298000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 85946 297200 86002 298000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 93674 297200 93730 298000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 101310 297200 101366 298000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 109038 297200 109094 298000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 116766 297200 116822 298000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 124494 297200 124550 298000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 132222 297200 132278 298000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 139858 297200 139914 298000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 147586 297200 147642 298000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 8850 297200 8906 298000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 155314 297200 155370 298000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 163042 297200 163098 298000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 170678 297200 170734 298000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 178406 297200 178462 298000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 186134 297200 186190 298000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 193862 297200 193918 298000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 201498 297200 201554 298000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 209226 297200 209282 298000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 216954 297200 217010 298000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 224682 297200 224738 298000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 16578 297200 16634 298000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 232410 297200 232466 298000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 240046 297200 240102 298000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 247774 297200 247830 298000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 255502 297200 255558 298000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 263230 297200 263286 298000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 270866 297200 270922 298000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 278594 297200 278650 298000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 286322 297200 286378 298000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 24306 297200 24362 298000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 32034 297200 32090 298000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 39670 297200 39726 298000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 47398 297200 47454 298000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 55126 297200 55182 298000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 62854 297200 62910 298000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 70490 297200 70546 298000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3698 297200 3754 298000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 80794 297200 80850 298000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 88522 297200 88578 298000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 96250 297200 96306 298000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 103886 297200 103942 298000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 111614 297200 111670 298000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 119342 297200 119398 298000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 127070 297200 127126 298000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 134706 297200 134762 298000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 142434 297200 142490 298000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 150162 297200 150218 298000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 11426 297200 11482 298000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 157890 297200 157946 298000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 165618 297200 165674 298000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 173254 297200 173310 298000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 180982 297200 181038 298000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 188710 297200 188766 298000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 196438 297200 196494 298000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 204074 297200 204130 298000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 211802 297200 211858 298000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 219530 297200 219586 298000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 227258 297200 227314 298000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 19154 297200 19210 298000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 234894 297200 234950 298000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 242622 297200 242678 298000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 250350 297200 250406 298000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 258078 297200 258134 298000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 265806 297200 265862 298000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 273442 297200 273498 298000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 281170 297200 281226 298000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 288898 297200 288954 298000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 26882 297200 26938 298000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 34518 297200 34574 298000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 42246 297200 42302 298000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 49974 297200 50030 298000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 57702 297200 57758 298000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 65430 297200 65486 298000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 73066 297200 73122 298000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 6274 297200 6330 298000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 83370 297200 83426 298000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 91098 297200 91154 298000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 98826 297200 98882 298000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 106462 297200 106518 298000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 114190 297200 114246 298000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 121918 297200 121974 298000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 129646 297200 129702 298000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 137282 297200 137338 298000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 145010 297200 145066 298000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 152738 297200 152794 298000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 14002 297200 14058 298000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 160466 297200 160522 298000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 168102 297200 168158 298000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 175830 297200 175886 298000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 183558 297200 183614 298000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 191286 297200 191342 298000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 199014 297200 199070 298000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 206650 297200 206706 298000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 214378 297200 214434 298000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 222106 297200 222162 298000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 229834 297200 229890 298000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 21730 297200 21786 298000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 237470 297200 237526 298000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 245198 297200 245254 298000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 252926 297200 252982 298000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 260654 297200 260710 298000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 268290 297200 268346 298000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 276018 297200 276074 298000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 283746 297200 283802 298000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 291474 297200 291530 298000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 29458 297200 29514 298000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 37094 297200 37150 298000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 44822 297200 44878 298000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 52550 297200 52606 298000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 60278 297200 60334 298000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 67914 297200 67970 298000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 75642 297200 75698 298000 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 0 148928 800 149048 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 294050 297200 294106 298000 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 296626 297200 296682 298000 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 64602 0 64658 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 246670 0 246726 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 248510 0 248566 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 250258 0 250314 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 252098 0 252154 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 253938 0 253994 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 255778 0 255834 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 257618 0 257674 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 259366 0 259422 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 261206 0 261262 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 263046 0 263102 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 264886 0 264942 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 266634 0 266690 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 268474 0 268530 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 270314 0 270370 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 272154 0 272210 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 273994 0 274050 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 275742 0 275798 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 277582 0 277638 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 279422 0 279478 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 281262 0 281318 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 283102 0 283158 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 284850 0 284906 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 286690 0 286746 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 288530 0 288586 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 290370 0 290426 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 292210 0 292266 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 293958 0 294014 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 295798 0 295854 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 120998 0 121054 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 128266 0 128322 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 131946 0 132002 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 135626 0 135682 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 142894 0 142950 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 146482 0 146538 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 157430 0 157486 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 159270 0 159326 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 161110 0 161166 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 162858 0 162914 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 166538 0 166594 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 168378 0 168434 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 171966 0 172022 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 173806 0 173862 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 175646 0 175702 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 177486 0 177542 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 179326 0 179382 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 181074 0 181130 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 182914 0 182970 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 184754 0 184810 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 186594 0 186650 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 188342 0 188398 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 190182 0 190238 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 192022 0 192078 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 195702 0 195758 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 197450 0 197506 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 199290 0 199346 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 201130 0 201186 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 202970 0 203026 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 204810 0 204866 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 206558 0 206614 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 208398 0 208454 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 210238 0 210294 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 212078 0 212134 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 213918 0 213974 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 215666 0 215722 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 217506 0 217562 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 219346 0 219402 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 221186 0 221242 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 223026 0 223082 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 224774 0 224830 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 226614 0 226670 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 228454 0 228510 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 230294 0 230350 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 232042 0 232098 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 233882 0 233938 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 235722 0 235778 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 237562 0 237618 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 239402 0 239458 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 241150 0 241206 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 242990 0 243046 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 244830 0 244886 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 247222 0 247278 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 249062 0 249118 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 250902 0 250958 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 252742 0 252798 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 254582 0 254638 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 256330 0 256386 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 258170 0 258226 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 260010 0 260066 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 261850 0 261906 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 263598 0 263654 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 83370 0 83426 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 265438 0 265494 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 267278 0 267334 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 269118 0 269174 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 270958 0 271014 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 272706 0 272762 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 274546 0 274602 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 276386 0 276442 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 278226 0 278282 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 280066 0 280122 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 281814 0 281870 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 283654 0 283710 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 285494 0 285550 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 287334 0 287390 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 289174 0 289230 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 290922 0 290978 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 292762 0 292818 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 294602 0 294658 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 296442 0 296498 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 87050 0 87106 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 96158 0 96214 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 97998 0 98054 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 99746 0 99802 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 101586 0 101642 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 103426 0 103482 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 105266 0 105322 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 110694 0 110750 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 112534 0 112590 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 116122 0 116178 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 117962 0 118018 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 121642 0 121698 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 123482 0 123538 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 125230 0 125286 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 127070 0 127126 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 128910 0 128966 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 132590 0 132646 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 134338 0 134394 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 136178 0 136234 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 70674 0 70730 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 138018 0 138074 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 139858 0 139914 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 141698 0 141754 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 143446 0 143502 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 145286 0 145342 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 147126 0 147182 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 148966 0 149022 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 152554 0 152610 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 154394 0 154450 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 72514 0 72570 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 156234 0 156290 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 158074 0 158130 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 159822 0 159878 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 161662 0 161718 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 163502 0 163558 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 165342 0 165398 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 167182 0 167238 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 168930 0 168986 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 170770 0 170826 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 172610 0 172666 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 174450 0 174506 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 176290 0 176346 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 178038 0 178094 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 179878 0 179934 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 181718 0 181774 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 183558 0 183614 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 185398 0 185454 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 187146 0 187202 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 188986 0 189042 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 190826 0 190882 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 192666 0 192722 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 194414 0 194470 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 196254 0 196310 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 198094 0 198150 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 199934 0 199990 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 201774 0 201830 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 203522 0 203578 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 205362 0 205418 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 207202 0 207258 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 209042 0 209098 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 210882 0 210938 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 212630 0 212686 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 214470 0 214526 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 216310 0 216366 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 218150 0 218206 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 219990 0 220046 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 221738 0 221794 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 223578 0 223634 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 225418 0 225474 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 227258 0 227314 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 79782 0 79838 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 229006 0 229062 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 230846 0 230902 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 232686 0 232742 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 234526 0 234582 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 236366 0 236422 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 238114 0 238170 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 239954 0 240010 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 241794 0 241850 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 243634 0 243690 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 245474 0 245530 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 247866 0 247922 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 249706 0 249762 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 251546 0 251602 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 253294 0 253350 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 255134 0 255190 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 256974 0 257030 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 258814 0 258870 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 260654 0 260710 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 262402 0 262458 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 264242 0 264298 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 266082 0 266138 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 267922 0 267978 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 269670 0 269726 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 271510 0 271566 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 273350 0 273406 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 275190 0 275246 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 277030 0 277086 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 278778 0 278834 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 280618 0 280674 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 282458 0 282514 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 284298 0 284354 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 286138 0 286194 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 287886 0 287942 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 289726 0 289782 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 291566 0 291622 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 293406 0 293462 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 295246 0 295302 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 296994 0 297050 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 116766 0 116822 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 122194 0 122250 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 124034 0 124090 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 125874 0 125930 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 129554 0 129610 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 134982 0 135038 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 138662 0 138718 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 144090 0 144146 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 151358 0 151414 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 156786 0 156842 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 158626 0 158682 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 160466 0 160522 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 162306 0 162362 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 164146 0 164202 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 165894 0 165950 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 167734 0 167790 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 169574 0 169630 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 171414 0 171470 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 173254 0 173310 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 175002 0 175058 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 180522 0 180578 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 182362 0 182418 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 184110 0 184166 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 185950 0 186006 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 187790 0 187846 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 189630 0 189686 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 191378 0 191434 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 193218 0 193274 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 195058 0 195114 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 196898 0 196954 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 198738 0 198794 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 200486 0 200542 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 202326 0 202382 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 204166 0 204222 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 206006 0 206062 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 207846 0 207902 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 209594 0 209650 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 211434 0 211490 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 213274 0 213330 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 215114 0 215170 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 216954 0 217010 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 218702 0 218758 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 220542 0 220598 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 222382 0 222438 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 224222 0 224278 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 225970 0 226026 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 227810 0 227866 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 229650 0 229706 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 231490 0 231546 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 233330 0 233386 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 235078 0 235134 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 236918 0 236974 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 238758 0 238814 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 240598 0 240654 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 242438 0 242494 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 244186 0 244242 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 246026 0 246082 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 297638 0 297694 800 6 user_clk
port 502 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 503 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 504 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_ack_o
port 505 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 wbs_adr_i[0]
port 506 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[10]
port 507 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_adr_i[11]
port 508 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_adr_i[12]
port 509 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_adr_i[13]
port 510 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_adr_i[14]
port 511 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_adr_i[15]
port 512 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_adr_i[16]
port 513 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_adr_i[17]
port 514 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wbs_adr_i[18]
port 515 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 wbs_adr_i[19]
port 516 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_adr_i[1]
port 517 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 wbs_adr_i[20]
port 518 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 wbs_adr_i[21]
port 519 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 wbs_adr_i[22]
port 520 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 wbs_adr_i[23]
port 521 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 wbs_adr_i[24]
port 522 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 wbs_adr_i[25]
port 523 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 wbs_adr_i[26]
port 524 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 wbs_adr_i[27]
port 525 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 wbs_adr_i[28]
port 526 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 wbs_adr_i[29]
port 527 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[2]
port 528 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 wbs_adr_i[30]
port 529 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 wbs_adr_i[31]
port 530 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_adr_i[3]
port 531 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_adr_i[4]
port 532 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_adr_i[5]
port 533 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_adr_i[6]
port 534 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_adr_i[7]
port 535 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[8]
port 536 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_adr_i[9]
port 537 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_cyc_i
port 538 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_dat_i[0]
port 539 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_i[10]
port 540 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_i[11]
port 541 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_i[12]
port 542 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 wbs_dat_i[13]
port 543 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_dat_i[14]
port 544 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 wbs_dat_i[15]
port 545 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_i[16]
port 546 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_i[17]
port 547 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 wbs_dat_i[18]
port 548 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 wbs_dat_i[19]
port 549 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_i[1]
port 550 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 wbs_dat_i[20]
port 551 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 wbs_dat_i[21]
port 552 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 wbs_dat_i[22]
port 553 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 wbs_dat_i[23]
port 554 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 wbs_dat_i[24]
port 555 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 wbs_dat_i[25]
port 556 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 wbs_dat_i[26]
port 557 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 wbs_dat_i[27]
port 558 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 wbs_dat_i[28]
port 559 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 wbs_dat_i[29]
port 560 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_i[2]
port 561 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 wbs_dat_i[30]
port 562 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 wbs_dat_i[31]
port 563 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_i[3]
port 564 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_i[4]
port 565 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_dat_i[5]
port 566 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_dat_i[6]
port 567 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_i[7]
port 568 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_i[8]
port 569 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_i[9]
port 570 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_o[0]
port 571 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_o[10]
port 572 nsew signal output
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_o[11]
port 573 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_o[12]
port 574 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_o[13]
port 575 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 wbs_dat_o[14]
port 576 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_o[15]
port 577 nsew signal output
rlabel metal2 s 36634 0 36690 800 6 wbs_dat_o[16]
port 578 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 wbs_dat_o[17]
port 579 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 wbs_dat_o[18]
port 580 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 wbs_dat_o[19]
port 581 nsew signal output
rlabel metal2 s 7562 0 7618 800 6 wbs_dat_o[1]
port 582 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 wbs_dat_o[20]
port 583 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 wbs_dat_o[21]
port 584 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 wbs_dat_o[22]
port 585 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 wbs_dat_o[23]
port 586 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 wbs_dat_o[24]
port 587 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 wbs_dat_o[25]
port 588 nsew signal output
rlabel metal2 s 54850 0 54906 800 6 wbs_dat_o[26]
port 589 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 wbs_dat_o[27]
port 590 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 wbs_dat_o[28]
port 591 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 wbs_dat_o[29]
port 592 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[2]
port 593 nsew signal output
rlabel metal2 s 62118 0 62174 800 6 wbs_dat_o[30]
port 594 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 wbs_dat_o[31]
port 595 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_o[3]
port 596 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[4]
port 597 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_o[5]
port 598 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_o[6]
port 599 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 wbs_dat_o[7]
port 600 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_o[8]
port 601 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_o[9]
port 602 nsew signal output
rlabel metal2 s 5722 0 5778 800 6 wbs_sel_i[0]
port 603 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_sel_i[1]
port 604 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_sel_i[2]
port 605 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_sel_i[3]
port 606 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_stb_i
port 607 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_we_i
port 608 nsew signal input
rlabel metal4 s 280688 2128 281008 295440 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 295440 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 295440 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 295440 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 295440 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 295440 6 vccd1
port 614 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 295440 6 vccd1
port 615 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 295440 6 vccd1
port 616 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 295440 6 vccd1
port 617 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 295440 6 vccd1
port 618 nsew power bidirectional
rlabel metal4 s 296048 2128 296368 295440 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 295440 6 vssd1
port 620 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 295440 6 vssd1
port 621 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 295440 6 vssd1
port 622 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 295440 6 vssd1
port 623 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 295440 6 vssd1
port 624 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 295440 6 vssd1
port 625 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 295440 6 vssd1
port 626 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 295440 6 vssd1
port 627 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 295440 6 vssd1
port 628 nsew ground bidirectional
rlabel metal4 s 281348 2176 281668 295392 6 vccd2
port 629 nsew power bidirectional
rlabel metal4 s 250628 2176 250948 295392 6 vccd2
port 630 nsew power bidirectional
rlabel metal4 s 219908 2176 220228 295392 6 vccd2
port 631 nsew power bidirectional
rlabel metal4 s 189188 2176 189508 295392 6 vccd2
port 632 nsew power bidirectional
rlabel metal4 s 158468 2176 158788 295392 6 vccd2
port 633 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 295392 6 vccd2
port 634 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 295392 6 vccd2
port 635 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 295392 6 vccd2
port 636 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 295392 6 vccd2
port 637 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 295392 6 vccd2
port 638 nsew power bidirectional
rlabel metal4 s 265988 2176 266308 295392 6 vssd2
port 639 nsew ground bidirectional
rlabel metal4 s 235268 2176 235588 295392 6 vssd2
port 640 nsew ground bidirectional
rlabel metal4 s 204548 2176 204868 295392 6 vssd2
port 641 nsew ground bidirectional
rlabel metal4 s 173828 2176 174148 295392 6 vssd2
port 642 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 295392 6 vssd2
port 643 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 295392 6 vssd2
port 644 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 295392 6 vssd2
port 645 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 295392 6 vssd2
port 646 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 295392 6 vssd2
port 647 nsew ground bidirectional
rlabel metal4 s 282008 2176 282328 295392 6 vdda1
port 648 nsew power bidirectional
rlabel metal4 s 251288 2176 251608 295392 6 vdda1
port 649 nsew power bidirectional
rlabel metal4 s 220568 2176 220888 295392 6 vdda1
port 650 nsew power bidirectional
rlabel metal4 s 189848 2176 190168 295392 6 vdda1
port 651 nsew power bidirectional
rlabel metal4 s 159128 2176 159448 295392 6 vdda1
port 652 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 295392 6 vdda1
port 653 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 295392 6 vdda1
port 654 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 295392 6 vdda1
port 655 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 295392 6 vdda1
port 656 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 295392 6 vdda1
port 657 nsew power bidirectional
rlabel metal4 s 266648 2176 266968 295392 6 vssa1
port 658 nsew ground bidirectional
rlabel metal4 s 235928 2176 236248 295392 6 vssa1
port 659 nsew ground bidirectional
rlabel metal4 s 205208 2176 205528 295392 6 vssa1
port 660 nsew ground bidirectional
rlabel metal4 s 174488 2176 174808 295392 6 vssa1
port 661 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 295392 6 vssa1
port 662 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 295392 6 vssa1
port 663 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 295392 6 vssa1
port 664 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 295392 6 vssa1
port 665 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 295392 6 vssa1
port 666 nsew ground bidirectional
rlabel metal4 s 282668 2176 282988 295392 6 vdda2
port 667 nsew power bidirectional
rlabel metal4 s 251948 2176 252268 295392 6 vdda2
port 668 nsew power bidirectional
rlabel metal4 s 221228 2176 221548 295392 6 vdda2
port 669 nsew power bidirectional
rlabel metal4 s 190508 2176 190828 295392 6 vdda2
port 670 nsew power bidirectional
rlabel metal4 s 159788 2176 160108 295392 6 vdda2
port 671 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 295392 6 vdda2
port 672 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 295392 6 vdda2
port 673 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 295392 6 vdda2
port 674 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 295392 6 vdda2
port 675 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 295392 6 vdda2
port 676 nsew power bidirectional
rlabel metal4 s 267308 2176 267628 295392 6 vssa2
port 677 nsew ground bidirectional
rlabel metal4 s 236588 2176 236908 295392 6 vssa2
port 678 nsew ground bidirectional
rlabel metal4 s 205868 2176 206188 295392 6 vssa2
port 679 nsew ground bidirectional
rlabel metal4 s 175148 2176 175468 295392 6 vssa2
port 680 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 295392 6 vssa2
port 681 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 295392 6 vssa2
port 682 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 295392 6 vssa2
port 683 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 295392 6 vssa2
port 684 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 295392 6 vssa2
port 685 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 298000 298000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 268376416
string GDS_START 834078
<< end >>

