`default_nettype none
//-----------------------------------------------------
// Project Name : a.out
// Function     : Main processor 
// Description  : This is the main processor
// Coder        : Jaquer AND VORIXO

//***Headers***
//***Module***
module decoder_output #(
        parameter integer WORD_SIZE = 32
    )
    (
        `ifdef USE_POWER_PINS
        inout vdda1,	// User area 1 3.3V supply
        inout vdda2,	// User area 2 3.3V supply
        inout vssa1,	// User area 1 analog ground
        inout vssa2,	// User area 2 analog ground
        inout vccd1,	// User area 1 1.8V supply
        inout vccd2,	// User area 2 1.8v supply
        inout vssd1,	// User area 1 digital ground
        inout vssd2,	// User area 2 digital ground
        `endif
        input  [1 : 0] operation_result_i ,
        input  [WORD_SIZE - 1 : 0] store_data_i ,
        output [1 : 0] operation_result_o ,
        output [WORD_SIZE - 1 : 0] store_data_o 
    );

//***Internal logic generated by compiler***  
    

//***Dumped Internal logic***
    assign operation_result_o = operation_result_i;
    assign store_data_o = store_data_i;

    
//***Handcrafted Internal logic*** 
//TODO
endmodule
